package background is 

TYPE my_background is array(0 to 79, 0 to 79) of integer range 0 to 250;

CONSTANT BASE_R: my_background :=
((76,73,75,76,76,79,74,72,78,75,77,75,72,69,71,76,76,84,86,70,75,76,76,76,74,76,72,73,71,73,70,76,73,68,73,76,80,81,72,77,78,74,74,72,76,83,74,71,78,79,79,74,74,76,78,74,77,78,76,73,74,75,72,75,70,72,75,70,76,72,78,82,71,73,75,74,73,74,76,74),
(77,73,73,73,72,77,77,76,74,68,73,74,75,75,84,77,67,73,75,81,76,73,69,68,64,75,79,75,77,75,80,77,74,80,80,73,73,79,71,76,79,75,78,75,75,72,76,80,68,72,70,81,80,77,77,72,74,78,76,92,83,69,77,79,78,85,82,74,78,74,75,70,80,75,73,75,77,70,74,75),
(78,82,84,83,86,73,125,119,83,73,73,89,83,81,128,118,87,83,99,130,106,86,82,79,84,117,134,82,81,88,88,87,69,109,131,90,79,79,85,86,75,110,136,88,82,80,122,127,81,80,86,134,124,72,80,83,92,82,74,126,118,75,81,79,89,82,74,124,124,82,81,87,134,111,84,86,81,72,75,77),
(68,80,88,79,78,70,129,119,83,75,69,89,77,74,132,121,81,74,85,138,112,78,81,80,82,116,134,83,84,89,77,78,65,116,132,83,81,72,86,86,64,109,138,85,70,72,127,135,88,81,84,134,121,69,89,86,88,75,71,134,117,91,79,68,82,72,68,133,127,77,69,82,141,119,80,79,70,69,74,76),
(84,85,84,91,82,76,120,107,76,87,82,82,77,77,122,119,82,87,96,131,110,81,84,84,78,114,119,74,72,87,93,91,72,104,125,96,86,80,83,80,68,105,130,89,84,91,116,122,89,80,84,123,109,82,85,80,94,86,77,117,121,101,90,80,78,84,92,130,113,83,87,95,123,113,85,81,86,87,79,74),
(125,83,76,131,108,77,98,88,74,116,123,82,84,84,93,90,70,103,127,85,79,78,77,79,72,84,88,86,78,76,117,121,84,91,98,120,146,129,86,76,87,90,94,79,98,134,101,86,76,78,80,81,101,128,88,77,127,113,82,88,90,100,126,128,86,95,99,96,97,78,114,125,95,85,75,76,95,133,98,78),
(138,90,83,141,113,80,84,84,77,126,133,86,85,81,79,75,68,130,138,76,87,72,80,82,74,75,81,82,79,83,128,126,82,83,81,125,145,142,100,86,81,78,78,78,96,141,95,76,75,82,85,73,105,149,94,75,137,107,69,76,90,94,124,134,75,94,105,86,76,58,117,124,80,78,76,77,93,146,104,79),
(136,101,91,129,98,76,83,83,82,121,126,81,73,80,94,93,67,121,137,79,80,66,74,79,81,86,88,80,71,78,115,119,83,79,80,135,136,126,99,89,83,84,94,79,88,131,95,78,73,81,87,80,103,144,91,74,125,104,76,83,92,107,126,124,82,100,103,84,81,62,128,138,76,75,78,82,94,129,102,81),
(110,107,103,85,74,71,81,75,77,79,82,78,90,93,101,90,91,95,106,107,94,87,85,91,134,93,71,83,74,67,76,86,74,77,84,92,92,84,68,71,82,86,98,89,82,86,82,81,75,82,84,76,72,83,75,76,86,78,74,85,95,165,119,103,68,105,174,120,116,90,98,108,97,75,73,83,74,74,74,72),
(111,110,103,79,80,82,85,81,87,79,77,72,74,77,111,99,86,92,109,103,93,70,73,90,143,105,80,85,78,80,81,87,73,70,71,118,98,77,71,73,82,101,118,90,76,88,87,83,76,81,89,80,78,88,73,76,84,84,70,72,94,164,132,98,75,112,148,103,105,91,97,105,90,76,82,90,82,79,86,78),
(127,122,116,87,86,86,76,86,97,90,82,77,82,77,114,100,69,114,134,122,117,89,90,98,125,98,80,87,85,84,85,88,87,79,68,115,92,86,87,91,96,106,101,91,79,76,77,84,82,85,83,82,83,92,75,77,91,87,84,75,97,159,111,92,91,113,150,120,109,68,112,112,79,81,92,78,70,83,89,93),
(153,141,145,126,117,87,85,90,91,93,83,98,114,112,131,99,68,150,193,192,151,88,123,123,76,97,104,83,89,111,106,104,101,95,89,111,93,74,91,101,96,108,100,77,78,87,84,69,80,81,79,107,100,83,81,87,92,100,110,94,95,161,111,92,110,127,162,156,136,61,156,181,87,82,102,81,88,138,103,89),
(161,152,150,133,127,115,93,92,121,79,70,110,107,103,108,102,70,160,198,192,154,104,139,124,80,104,104,83,83,110,102,114,112,93,87,112,99,63,117,115,99,118,114,70,70,81,81,68,87,78,82,100,105,74,71,93,119,114,101,78,97,174,93,67,107,133,162,142,135,63,150,197,81,90,111,81,89,145,114,103),
(155,140,139,145,113,118,89,94,124,97,85,110,116,114,103,108,75,156,191,191,157,118,126,109,80,107,116,84,94,118,116,111,116,97,79,108,110,78,97,111,115,117,115,80,75,66,74,89,93,81,87,102,101,78,84,90,118,112,104,94,100,141,99,80,110,126,154,138,138,74,151,188,67,92,127,83,90,121,118,120),
(130,96,89,90,130,154,70,93,161,119,114,163,152,156,148,133,101,129,163,190,168,152,80,89,99,150,153,98,123,161,147,150,155,105,70,106,109,120,76,102,159,148,148,114,105,102,119,99,71,86,114,170,139,84,80,84,143,154,164,115,102,78,111,118,175,162,152,92,71,101,132,147,70,107,169,120,96,81,127,160),
(140,94,77,117,141,160,81,101,159,118,109,164,161,165,142,118,104,132,163,200,184,148,92,79,105,135,155,110,124,157,154,158,165,109,69,108,110,111,83,93,158,154,155,110,103,66,93,115,73,92,110,154,134,62,78,89,153,152,150,112,96,71,101,118,151,155,156,106,100,115,145,148,76,110,159,117,99,83,134,165),
(133,107,89,100,126,152,83,101,141,130,125,159,154,156,123,119,112,130,150,169,173,149,101,94,115,145,151,130,131,147,152,155,136,98,98,116,125,112,93,108,163,157,158,121,98,80,99,119,78,105,125,148,134,88,88,100,139,157,142,123,113,87,98,101,160,159,154,93,96,117,140,149,84,110,177,131,100,71,131,162),
(163,119,98,87,125,155,117,106,78,124,145,159,155,156,88,98,167,93,73,132,149,155,102,112,160,160,155,152,158,159,142,131,88,98,103,152,159,162,104,111,155,149,152,166,123,63,127,140,78,122,153,161,142,103,115,100,88,109,155,157,136,109,87,90,158,162,157,105,105,148,152,147,146,136,137,144,138,72,128,162),
(155,124,111,63,110,158,116,102,53,124,158,154,156,154,88,96,171,107,88,145,137,158,120,127,159,157,158,152,151,157,165,136,67,106,125,154,146,156,125,119,148,149,147,163,130,64,114,128,71,120,158,152,132,98,117,108,65,102,167,145,141,119,82,85,153,161,162,121,118,159,155,147,136,150,156,160,131,66,124,162),
(142,122,106,79,127,158,96,97,101,143,163,151,153,154,93,96,142,97,78,142,145,152,127,125,149,151,160,154,147,149,154,131,81,101,119,154,142,144,124,130,160,155,145,153,126,84,121,137,82,121,160,165,158,118,116,113,85,124,163,142,136,103,98,111,154,154,155,118,125,162,149,159,121,142,153,166,129,78,132,165),
(160,168,146,103,139,167,168,149,102,133,151,151,150,154,115,103,80,105,126,135,148,153,149,149,148,154,160,148,161,163,92,73,118,138,158,157,151,160,184,192,199,173,144,164,127,94,151,142,64,115,158,151,165,158,160,142,115,128,160,157,149,168,115,98,153,155,143,153,153,149,152,150,100,121,129,150,154,100,136,157),
(154,155,146,104,131,152,150,142,109,130,154,153,152,148,110,93,82,83,115,161,152,150,154,155,155,156,158,152,154,159,79,77,89,136,159,152,159,158,181,193,192,169,154,163,137,111,146,131,71,113,155,149,153,150,158,147,103,120,159,158,156,156,131,113,149,154,148,156,152,152,154,152,114,112,132,152,148,104,143,160),
(143,142,143,118,139,155,153,147,137,158,162,150,155,153,127,110,98,111,118,146,148,154,154,152,157,157,155,148,144,157,101,98,131,150,158,155,154,151,176,185,182,167,154,159,144,117,150,138,91,126,157,148,157,164,146,143,119,134,153,155,154,151,138,123,146,159,166,163,154,152,156,145,121,119,135,131,133,130,154,157),
(139,137,143,147,155,158,143,165,190,193,184,154,153,149,156,137,94,146,150,108,129,156,155,154,156,154,155,155,153,166,107,119,204,193,181,155,154,151,156,150,152,155,153,150,149,141,160,144,88,134,160,146,165,190,156,150,150,153,154,156,153,152,151,148,148,172,197,192,177,152,153,152,159,125,112,82,99,202,163,147),
(132,131,137,153,153,154,149,167,201,193,188,155,149,143,158,147,109,153,150,102,133,158,150,151,151,149,153,154,151,163,115,128,205,191,194,153,151,149,147,151,155,159,157,150,155,149,155,158,101,136,157,148,168,198,164,147,154,157,154,151,152,152,158,164,152,173,187,192,185,150,155,152,154,144,89,80,101,202,163,150),
(133,132,140,151,155,151,157,163,181,179,183,157,156,156,161,148,119,131,154,109,136,160,151,154,154,152,157,158,153,152,133,128,199,193,177,156,154,154,154,156,145,139,138,144,150,156,142,138,108,132,155,151,166,181,168,158,154,155,154,152,153,153,152,148,145,158,172,193,187,148,155,149,148,149,138,81,94,199,169,150),
(136,139,141,145,153,155,193,184,149,149,152,148,174,199,192,192,193,162,151,111,131,156,151,160,189,197,184,160,149,150,181,195,193,164,151,153,155,160,153,144,115,106,106,107,127,152,115,107,107,130,154,157,147,146,178,192,190,171,151,156,155,152,154,145,139,133,134,176,185,153,155,145,142,172,198,128,134,206,168,151),
(133,136,135,149,151,152,186,181,155,153,155,152,170,199,186,187,196,174,147,110,134,155,152,161,187,192,190,150,153,152,183,197,191,167,147,148,153,156,152,142,107,107,109,106,128,158,113,103,106,135,157,149,154,149,176,195,198,175,151,153,155,150,155,156,141,131,133,182,189,143,154,154,150,168,193,114,132,201,168,151),
(138,140,141,157,150,143,170,166,151,153,153,154,170,193,177,173,173,159,145,107,127,139,150,165,180,182,184,164,165,154,167,167,177,160,144,146,156,154,155,143,122,116,113,125,130,151,142,137,121,132,142,155,159,155,171,180,181,164,155,150,153,153,143,135,134,141,145,181,174,136,154,157,155,166,190,127,129,178,158,146),
(153,154,150,157,148,139,147,146,151,154,154,150,171,189,152,144,142,147,148,106,110,112,139,151,155,155,157,190,176,151,118,130,161,139,141,135,144,154,153,149,152,126,110,149,152,151,185,187,156,126,108,150,157,158,156,154,154,154,156,150,152,155,132,106,106,130,140,158,154,142,153,160,155,148,152,143,140,147,147,148),
(157,156,152,156,146,133,129,136,154,154,153,147,173,190,140,133,134,146,152,109,108,110,141,153,150,151,156,202,176,148,112,118,163,135,133,129,141,153,152,151,157,129,108,143,151,147,185,188,162,131,102,151,160,159,155,150,151,152,154,152,153,156,130,106,107,138,147,153,146,139,142,151,152,155,150,143,129,127,146,155),
(151,152,149,157,144,128,130,139,153,153,153,150,169,181,141,135,135,149,155,126,121,125,144,159,155,153,154,178,162,137,131,131,152,158,150,134,145,149,151,151,154,134,120,149,151,152,183,186,154,134,118,139,140,136,149,152,152,153,154,154,155,154,138,123,109,132,154,156,145,141,140,141,136,142,154,153,139,127,148,156),
(147,153,154,159,145,134,139,143,151,153,149,146,151,143,141,140,134,144,157,157,156,160,156,153,154,154,151,154,132,101,175,190,148,156,149,129,140,151,153,155,159,156,146,155,155,157,179,184,155,154,156,112,107,104,137,151,150,153,156,154,157,148,152,150,114,127,150,151,154,154,145,135,99,130,151,148,142,133,149,152),
(152,150,152,156,142,140,141,146,155,157,150,149,156,147,140,137,134,147,157,153,149,151,153,154,154,154,151,157,137,110,172,182,148,156,148,141,144,157,155,153,154,152,146,154,154,153,179,191,154,150,151,115,114,111,138,157,158,150,154,153,151,149,153,148,106,130,152,151,154,152,141,134,108,130,153,151,146,138,150,154),
(156,144,140,152,134,125,141,145,152,157,152,141,142,139,146,146,146,149,155,152,151,151,152,153,153,153,151,156,136,108,169,179,149,153,149,149,141,131,147,144,146,150,150,154,154,153,182,190,167,156,146,126,121,111,129,141,157,150,153,148,145,151,154,151,127,134,139,152,154,147,131,128,113,132,157,151,150,145,151,154),
(153,128,118,155,130,106,139,149,153,155,145,115,107,110,145,155,155,151,154,151,153,154,152,153,153,153,151,156,137,104,148,160,150,156,153,154,139,102,135,137,138,148,153,153,153,153,179,190,191,172,147,152,137,108,114,118,151,151,152,142,141,152,152,153,153,135,114,145,151,146,118,110,106,132,159,149,153,152,153,155),
(162,121,105,168,130,105,156,160,154,156,147,116,107,113,147,154,155,151,153,150,153,154,149,150,149,151,151,156,137,102,140,153,154,154,152,157,139,101,131,136,135,147,155,153,153,156,188,198,199,181,148,162,136,103,105,113,156,154,152,137,139,152,151,153,158,131,101,146,146,141,116,107,104,126,156,148,154,155,154,155),
(144,127,127,145,131,127,147,155,152,153,148,131,115,108,147,155,151,149,153,153,156,152,163,162,164,163,154,159,135,104,150,158,152,150,151,154,137,106,131,133,134,146,159,155,146,135,158,169,180,166,152,153,137,124,117,124,153,154,152,134,142,145,155,152,150,135,119,150,145,137,128,127,129,130,151,151,151,153,153,153),
(102,142,156,103,134,160,153,154,155,151,154,159,129,106,147,154,152,151,153,150,153,155,190,194,197,170,152,159,137,105,147,161,150,153,150,154,138,105,131,135,136,144,154,157,137,105,106,110,150,151,154,150,151,153,154,152,151,152,149,128,134,139,145,148,154,153,155,149,146,148,154,158,156,153,154,153,153,153,153,153),
(107,142,148,105,133,163,158,152,157,151,150,157,128,107,148,152,154,156,153,153,152,157,193,195,193,159,148,158,138,109,140,156,154,152,149,151,137,101,133,138,139,144,150,156,141,105,115,124,150,155,153,150,152,151,151,153,150,146,148,141,138,133,142,152,156,155,149,148,157,160,154,151,157,155,153,149,151,153,153,153),
(127,145,152,127,142,158,151,147,154,154,152,158,134,110,147,153,154,151,153,174,161,155,169,175,187,174,167,157,142,129,146,152,169,169,173,155,134,103,128,134,143,146,151,157,137,108,123,132,151,152,151,155,152,155,157,154,147,147,152,163,162,136,152,151,134,147,152,154,150,149,149,148,158,150,151,145,151,153,153,153),
(151,153,154,145,153,155,140,143,152,154,153,160,131,110,148,155,152,151,154,189,174,152,154,161,192,191,184,155,151,149,154,163,193,192,189,156,135,108,103,113,146,148,153,156,139,115,143,156,155,152,152,154,153,153,153,153,153,151,153,180,171,129,150,148,111,136,153,156,152,149,152,149,154,144,137,134,143,152,153,153),
(156,153,153,157,155,150,138,137,155,153,151,153,130,107,149,154,154,155,150,191,176,150,152,165,200,195,188,153,155,156,152,167,198,188,184,158,139,105,100,118,154,160,156,155,136,109,145,153,142,154,155,155,154,155,154,152,157,151,156,192,171,131,147,152,108,132,153,154,152,153,156,151,150,148,136,126,140,148,153,152),
(153,153,152,151,152,149,144,140,149,148,154,168,147,122,150,156,154,154,164,194,174,152,153,158,171,180,175,157,157,156,152,158,177,180,187,160,145,122,123,134,153,159,150,157,136,122,145,146,141,148,146,152,150,137,151,152,152,152,155,189,182,157,154,150,110,132,155,152,149,152,156,149,154,150,149,144,148,143,152,158),
(153,153,152,152,153,153,153,147,136,144,157,195,176,150,154,155,156,177,194,197,174,154,155,155,149,147,148,156,155,155,154,152,145,178,196,156,152,154,153,152,151,153,146,152,155,151,140,134,142,135,136,150,138,106,142,154,150,153,153,189,198,188,165,145,111,131,155,152,153,153,157,147,152,150,152,155,143,133,145,159),
(153,153,153,153,155,154,158,150,129,146,161,192,172,150,153,149,150,175,190,196,173,153,157,154,157,157,156,154,149,156,153,154,157,177,183,151,147,149,151,149,152,152,158,154,156,155,136,126,133,126,130,150,135,105,145,158,156,152,156,189,198,195,167,139,110,130,156,152,156,152,151,149,150,150,155,160,147,134,142,154),
(152,153,154,153,152,151,156,148,131,146,163,194,176,152,154,147,128,173,192,176,164,154,156,154,153,145,137,137,144,157,153,153,150,176,193,173,161,154,157,152,147,145,157,149,152,161,152,144,140,150,150,156,145,125,127,135,152,150,155,169,173,179,149,124,108,132,157,151,161,173,169,171,171,161,151,154,151,145,147,156),
(152,153,154,154,154,151,152,148,134,145,162,191,174,149,152,144,106,166,191,155,155,153,149,151,157,129,107,109,132,158,152,152,154,174,195,191,173,154,156,150,134,142,153,148,155,156,156,151,137,147,150,150,154,153,117,121,154,150,151,150,147,154,126,113,107,130,154,151,165,193,189,191,196,178,154,156,159,148,147,152),
(153,153,153,153,155,155,149,150,143,147,156,190,171,146,153,138,102,170,200,157,158,154,149,154,156,127,103,106,125,159,154,154,152,178,194,193,180,152,152,149,132,147,158,147,148,151,153,148,137,138,148,152,157,158,122,116,152,151,152,152,156,152,126,107,108,131,155,149,161,191,189,187,195,180,150,153,152,155,155,154),
(153,153,153,154,154,157,142,146,154,148,158,184,177,167,159,142,112,138,153,133,140,153,160,153,134,116,106,132,140,156,154,154,152,169,173,173,168,153,152,150,142,144,147,150,155,152,151,154,146,147,152,157,150,132,126,130,152,152,154,153,155,152,138,128,128,143,154,151,158,174,185,184,178,166,149,154,153,154,154,154),
(153,153,153,154,154,154,134,137,151,152,161,190,197,189,161,140,109,109,98,103,129,156,156,141,103,104,110,153,158,152,148,154,154,150,151,150,152,152,153,150,134,134,138,151,155,151,154,155,147,148,153,160,135,101,138,156,153,152,154,154,154,151,152,157,151,153,154,153,154,152,182,190,153,150,152,153,153,154,154,154),
(153,153,153,155,154,152,137,140,150,155,160,189,187,186,162,138,108,108,105,103,126,154,155,145,107,107,112,150,160,152,150,152,155,152,157,156,158,154,152,149,130,134,141,151,155,150,158,154,151,151,152,158,137,106,142,151,151,155,153,154,156,152,151,151,150,152,154,154,155,150,178,192,154,155,155,153,153,154,154,154),
(153,153,153,155,154,152,147,153,156,155,154,174,184,193,159,144,134,127,131,134,145,153,151,143,137,138,135,147,152,155,158,152,152,157,155,154,154,154,153,150,137,144,148,132,133,128,142,151,159,156,151,151,148,139,148,156,152,156,151,154,153,153,154,154,156,155,154,154,155,153,165,173,158,154,153,153,153,154,154,154),
(154,153,152,150,152,152,154,156,151,154,153,146,170,197,155,154,157,154,158,154,154,151,150,156,154,154,152,152,147,151,156,154,154,159,153,151,154,156,152,145,134,145,148,113,106,116,138,148,153,159,152,153,153,153,153,154,155,152,150,161,157,154,155,154,154,153,154,153,151,153,154,152,152,149,152,149,157,157,154,153),
(153,153,152,150,154,157,149,150,154,153,154,146,168,194,154,151,153,153,154,154,155,150,150,157,154,152,154,154,152,152,154,157,150,152,154,152,155,153,145,143,142,149,154,113,112,116,139,152,151,160,152,154,156,154,156,155,153,153,151,155,156,153,153,154,154,154,154,153,151,153,154,153,152,150,153,146,156,155,154,152),
(153,152,151,154,145,131,143,153,154,153,154,149,172,194,155,151,153,154,153,154,157,152,134,139,154,155,157,156,154,154,136,135,150,154,154,152,154,150,144,141,145,148,154,135,122,106,142,147,129,146,153,157,159,158,155,154,156,143,129,152,154,149,151,153,153,153,153,152,151,153,154,153,152,151,154,132,137,156,153,151),
(152,151,150,155,130,105,143,155,151,153,154,152,174,193,159,156,157,155,153,154,156,154,119,119,151,156,155,153,151,152,117,114,152,158,153,152,153,150,143,142,144,147,152,161,139,104,144,143,108,131,155,157,157,157,152,151,158,131,106,148,153,149,150,152,152,153,152,150,151,153,154,153,153,152,154,119,117,157,153,150),
(152,152,153,156,127,113,146,148,151,152,155,150,169,188,158,154,152,153,154,154,154,154,121,120,154,156,153,150,151,155,117,122,151,151,154,152,153,153,137,146,151,155,153,151,142,107,140,152,112,133,158,157,154,153,155,155,157,133,114,144,154,150,151,152,152,153,152,151,152,153,154,153,153,153,155,123,120,155,152,150),
(152,143,137,134,124,108,149,153,153,153,154,149,162,174,139,138,150,155,156,154,156,154,111,114,162,144,147,159,147,133,110,117,156,152,153,153,153,152,147,145,133,145,153,153,150,129,149,149,103,131,162,141,153,159,141,136,139,118,108,136,148,154,150,152,153,153,149,145,145,153,153,154,153,154,157,113,112,156,150,148),
(160,123,108,109,109,110,136,137,150,154,153,153,156,147,110,123,156,155,155,154,155,152,117,121,163,142,138,150,131,107,111,116,139,139,153,153,153,152,148,136,108,134,157,155,155,151,153,145,107,137,160,138,141,151,122,111,114,112,106,134,148,154,153,152,152,155,152,118,121,153,152,149,156,153,152,119,117,154,143,140),
(156,117,102,112,111,105,129,137,152,153,153,151,155,149,107,122,162,157,153,155,152,155,117,117,152,140,138,150,126,106,108,111,133,141,154,153,153,156,154,140,106,138,164,156,152,149,153,150,106,130,153,137,142,148,116,109,113,104,102,133,144,151,154,152,153,153,152,119,122,151,157,156,155,152,154,119,118,153,137,130),
(152,139,130,131,129,133,143,147,160,152,153,153,156,148,111,116,131,129,131,153,152,153,137,138,150,142,146,155,144,129,128,135,143,152,158,152,153,151,154,142,102,120,135,129,139,151,153,153,132,144,148,142,149,154,136,131,132,130,129,140,145,148,154,152,152,153,153,115,112,132,130,131,150,154,152,137,138,162,151,143),
(153,157,160,154,153,157,152,155,155,153,153,151,155,152,116,107,104,104,112,152,153,149,156,153,154,150,155,154,155,154,156,154,152,156,154,153,153,149,156,143,110,106,104,106,125,157,157,154,153,153,153,152,155,153,156,157,152,160,161,151,153,150,156,152,152,154,152,117,107,112,105,111,143,153,148,154,156,151,149,154),
(150,152,154,157,156,148,153,159,152,153,153,152,155,148,118,113,108,111,115,153,151,151,154,152,153,152,154,154,149,156,151,149,156,157,153,153,153,151,156,142,112,110,109,112,124,156,153,154,154,151,153,151,154,150,151,157,155,149,155,160,153,152,156,152,153,154,152,117,107,109,109,118,146,150,147,150,155,149,150,157),
(152,153,154,157,154,150,149,152,156,135,131,154,154,154,141,125,103,128,135,151,165,172,155,154,155,135,129,154,158,156,152,151,150,154,154,128,138,156,154,151,138,118,107,132,139,156,168,169,152,156,151,128,136,157,153,152,158,160,150,149,155,154,137,136,151,153,155,140,126,104,124,138,152,157,172,160,154,154,137,125),
(152,153,153,145,151,154,151,154,154,121,115,151,152,155,155,137,109,140,156,152,172,192,158,149,159,123,115,147,151,144,151,154,150,156,147,113,126,155,152,156,153,126,113,149,155,154,182,186,150,154,153,114,126,152,156,150,147,153,152,156,156,157,124,111,150,153,151,152,143,108,137,162,151,167,196,162,153,154,128,108),
(152,154,152,150,154,154,149,146,151,122,118,148,154,152,151,141,108,133,149,145,170,202,159,150,159,122,110,146,151,151,153,155,146,149,145,115,126,153,153,151,151,130,110,141,150,145,187,192,151,154,153,110,122,152,154,158,155,149,154,153,148,151,126,114,153,155,152,152,140,105,130,149,147,171,197,166,151,151,127,109),
(151,154,150,124,141,158,173,173,179,138,132,154,153,152,150,152,138,162,174,174,171,165,153,152,156,125,113,151,145,123,147,165,174,176,172,129,140,155,152,151,151,148,141,170,173,174,169,162,151,154,152,114,124,154,157,152,129,135,156,174,176,175,148,131,151,155,153,155,150,129,156,178,181,173,169,155,154,154,128,107),
(153,154,150,107,132,157,189,194,198,166,154,156,151,156,157,153,150,178,195,197,174,151,155,151,157,124,112,154,143,103,139,164,195,194,194,157,156,154,151,158,155,152,153,189,194,197,162,154,152,154,152,112,123,156,157,141,110,128,157,191,199,200,171,153,149,153,154,152,155,152,179,195,197,175,152,151,154,156,130,109),
(153,158,151,114,132,157,186,187,192,168,151,156,154,155,154,150,152,175,190,188,174,154,149,150,157,121,111,150,136,108,139,162,191,186,191,158,153,155,154,155,152,150,155,183,189,187,166,153,148,154,151,110,120,152,153,143,114,129,157,183,189,189,163,152,151,156,154,153,149,151,180,191,198,177,144,153,154,155,126,107),
(153,144,129,109,126,157,171,176,188,163,155,157,152,150,154,156,153,167,175,193,175,152,149,157,178,131,111,152,136,106,141,162,173,180,185,156,158,155,151,151,155,155,155,171,178,195,164,152,148,165,172,114,122,153,136,128,111,133,157,166,181,191,166,152,154,154,156,156,156,149,165,177,196,178,151,152,157,179,136,107),
(154,119,102,108,134,154,150,167,194,159,149,153,154,151,151,155,150,151,160,193,175,151,150,163,197,138,109,151,135,109,149,160,150,178,190,150,152,152,155,150,153,154,150,152,169,195,164,151,149,176,190,117,122,155,116,106,105,134,155,146,156,194,167,152,153,153,152,151,158,157,152,154,195,178,146,151,163,198,141,106),
(156,119,108,101,125,155,145,170,199,164,149,153,153,153,156,158,156,158,159,190,175,151,149,160,196,135,108,150,134,108,140,152,147,183,193,155,151,153,154,154,157,158,157,156,167,193,164,151,148,173,189,114,121,156,123,107,104,132,159,153,165,200,172,150,156,157,155,154,155,158,155,154,189,180,152,152,161,195,141,108),
(152,141,140,132,143,158,155,161,171,163,150,159,143,125,127,127,128,129,136,189,176,150,151,165,198,137,110,150,146,135,151,156,155,165,171,159,151,160,135,126,128,126,130,127,150,194,164,150,151,176,191,115,120,155,147,136,132,138,158,154,156,169,160,151,154,138,128,128,123,126,128,136,189,179,150,151,163,199,146,106),
(156,159,156,156,155,154,157,149,146,153,154,159,127,100,110,111,111,103,117,194,180,151,148,159,198,138,111,149,155,154,154,156,155,147,147,154,155,156,111,101,109,108,109,98,139,199,167,151,147,172,193,117,121,154,151,148,152,153,153,152,153,150,153,153,157,128,103,107,102,102,102,113,197,180,148,153,161,199,138,101),
(152,151,150,153,153,152,151,152,150,151,156,155,136,114,114,114,113,102,121,189,168,149,153,164,197,140,113,146,153,153,155,153,151,152,150,152,156,154,124,112,110,110,110,96,140,197,156,151,154,174,192,120,127,152,154,154,153,155,152,152,155,156,158,154,157,136,113,111,112,111,106,120,186,176,154,153,163,196,140,106),
(154,153,154,155,155,153,153,146,125,140,152,153,142,133,134,134,134,136,138,160,152,147,154,159,175,147,134,152,153,150,154,153,154,139,126,146,152,152,137,131,134,134,135,130,139,164,147,150,154,164,173,136,141,155,156,154,154,151,148,156,145,129,146,156,154,149,136,154,161,169,150,135,152,154,155,153,159,173,150,132),
(150,150,151,151,152,150,155,142,105,136,149,152,146,149,154,153,153,168,149,125,142,150,151,150,151,150,151,153,151,150,154,151,156,128,109,144,149,152,145,150,155,154,158,166,146,136,145,151,150,151,150,151,153,157,153,150,155,157,153,158,141,107,137,156,152,156,152,186,193,194,172,149,132,140,153,153,151,151,158,157),
(153,159,157,150,149,148,158,143,114,137,153,153,150,152,153,153,153,150,153,139,137,153,155,156,154,150,155,153,151,155,154,151,158,131,116,145,153,151,150,150,147,146,151,159,149,134,141,156,154,157,151,151,156,154,157,155,154,156,155,154,139,109,135,155,152,148,150,181,189,198,166,145,144,148,153,154,153,151,152,152),
(150,137,125,128,141,151,159,144,143,148,153,151,152,152,153,153,154,148,148,149,149,157,154,156,155,150,152,152,148,129,144,157,156,141,145,149,153,150,151,161,179,177,180,157,146,142,153,156,154,157,153,149,152,148,129,128,125,135,154,154,144,138,148,153,152,166,177,192,185,163,156,147,147,148,153,154,154,154,150,155));

CONSTANT BASE_G: my_background :=
((177,169,168,171,168,172,176,174,177,173,175,171,172,176,173,174,175,180,171,165,173,174,173,176,175,172,174,178,175,175,172,174,173,178,176,174,170,174,174,175,176,174,178,178,177,172,176,176,170,173,176,176,175,173,172,174,173,177,176,170,171,167,176,176,173,174,178,175,174,179,176,172,178,173,171,174,175,170,176,178),
(178,177,183,181,173,173,175,178,180,173,176,181,178,173,179,176,173,181,172,175,176,177,176,177,175,173,172,174,176,172,178,178,176,179,176,179,176,175,177,178,176,171,174,173,177,174,174,174,177,180,174,174,173,175,178,180,179,182,172,179,173,174,173,168,175,174,163,174,174,174,177,173,175,174,174,172,175,170,174,174),
(176,195,212,208,194,170,216,217,198,182,181,206,188,169,212,216,205,210,212,221,210,201,203,201,205,217,217,172,183,204,203,198,169,194,222,205,195,177,195,197,172,201,226,200,208,209,216,211,207,206,200,220,207,171,190,204,209,191,166,204,218,205,187,175,201,188,172,214,216,200,210,211,217,209,204,204,195,178,176,171),
(166,193,216,205,189,170,221,220,206,182,175,210,185,165,216,221,204,204,202,228,219,198,208,206,204,216,221,174,194,219,206,194,165,204,226,197,192,170,201,206,166,201,230,209,211,208,222,222,210,210,206,225,209,167,200,210,207,183,166,220,224,211,190,177,213,195,177,216,220,209,211,210,226,218,208,217,200,174,174,175),
(182,194,202,208,194,183,216,215,206,186,182,204,191,181,217,222,200,204,210,224,211,200,211,210,197,211,219,179,182,201,205,202,179,204,226,206,188,176,201,204,178,203,221,197,203,205,215,218,199,206,213,223,207,180,190,200,209,194,184,217,205,179,182,181,207,187,154,211,214,195,205,205,219,213,197,210,204,184,179,179),
(223,188,178,220,211,199,212,206,205,214,217,209,205,203,205,201,170,207,230,205,188,172,195,200,177,196,207,203,194,178,214,218,200,201,205,219,220,217,211,204,200,201,201,175,192,218,205,198,174,191,206,204,206,229,190,183,219,207,199,212,172,80,177,214,209,152,82,192,200,173,210,214,207,188,176,196,208,212,203,200),
(226,184,173,224,215,207,207,210,202,214,217,204,206,200,209,204,169,212,226,209,194,161,198,200,172,191,205,206,195,172,218,221,208,207,209,226,224,225,211,204,199,213,214,175,190,225,206,197,173,190,207,205,210,222,182,178,228,212,199,214,170,55,183,233,221,147,61,194,213,166,203,231,214,184,172,198,210,227,214,205),
(210,181,171,227,210,199,208,215,205,218,217,204,215,225,190,188,181,199,206,183,185,185,213,196,174,192,205,207,189,166,216,223,204,201,207,200,211,225,203,199,215,200,189,179,196,229,215,202,174,192,208,201,208,223,177,175,232,221,200,217,169,70,169,219,212,140,76,169,199,180,185,206,207,192,173,202,214,222,210,201),
(79,75,95,202,188,178,206,205,200,204,206,174,180,200,89,103,210,120,65,74,125,169,190,208,222,188,177,207,198,170,202,195,170,178,174,74,124,212,180,184,213,125,80,197,207,199,206,203,176,194,206,175,179,215,183,174,202,183,172,208,179,106,82,77,170,148,93,77,105,212,119,82,204,200,166,200,198,174,174,176),
(81,76,96,211,188,167,201,208,205,212,204,177,197,219,96,106,225,122,70,70,125,182,196,207,222,191,172,205,196,170,203,199,171,176,167,73,132,217,178,186,223,124,68,201,214,208,211,198,175,196,205,177,186,211,186,177,206,192,173,211,176,102,84,82,178,146,106,82,111,222,115,77,207,200,171,208,208,180,176,171),
(82,77,99,216,183,158,199,201,184,198,191,163,177,189,85,118,220,129,81,91,119,161,200,213,219,178,166,202,189,164,187,181,156,173,181,76,134,214,160,157,192,126,78,195,204,209,201,191,172,194,215,157,172,208,184,184,185,179,157,204,176,110,104,107,162,145,114,86,103,219,120,100,203,181,153,194,197,184,166,153),
(105,104,123,228,147,89,206,181,89,154,167,87,84,90,70,108,178,151,133,150,122,89,204,217,181,115,93,207,160,76,88,96,92,159,204,71,113,181,116,85,93,86,84,170,185,213,177,183,196,200,205,93,125,211,202,190,103,93,88,185,184,96,151,164,81,96,117,99,115,179,153,144,183,141,88,155,185,223,147,87),
(108,108,122,240,143,54,197,166,60,151,176,78,76,77,70,99,181,160,142,153,113,63,200,213,176,102,87,219,150,64,81,70,65,164,212,81,113,189,84,67,76,77,84,167,192,213,186,180,207,211,208,76,115,212,210,184,72,61,81,202,192,92,159,171,76,91,107,105,131,177,159,146,178,127,65,156,191,231,128,62),
(107,121,133,216,145,74,197,169,66,141,160,86,79,85,91,107,161,150,136,152,123,65,200,211,164,100,90,202,147,72,89,77,75,155,197,81,107,171,108,88,78,81,93,150,181,218,176,164,204,196,185,93,122,210,212,190,83,82,89,175,173,119,160,152,77,101,110,122,128,163,145,138,183,133,75,142,176,235,134,67),
(135,189,182,63,94,113,171,164,111,80,77,109,106,109,216,188,69,104,115,148,130,108,166,146,75,99,103,76,86,117,107,121,115,149,183,79,80,66,186,194,112,116,113,74,116,212,101,82,178,129,63,97,128,167,190,196,117,113,104,71,112,227,108,70,105,104,107,196,183,65,105,121,178,155,94,83,95,210,148,107),
(135,192,193,67,85,115,167,152,107,81,76,101,101,103,206,186,62,101,109,145,126,102,178,152,70,101,106,74,91,108,104,105,99,147,175,77,79,74,183,193,102,105,109,67,116,228,106,78,185,125,74,111,132,181,207,198,108,111,111,71,109,229,115,67,110,109,100,200,177,67,93,119,166,146,105,72,94,219,143,100),
(136,174,175,102,107,111,153,151,137,91,101,111,108,111,210,178,69,117,128,145,126,101,142,132,81,100,110,94,99,115,109,117,129,146,147,94,85,80,163,165,112,108,108,79,123,208,124,101,194,128,74,104,126,156,184,180,125,112,119,83,119,198,125,104,105,108,107,171,162,84,94,117,186,153,99,87,110,218,142,99),
(108,93,98,167,139,107,85,113,218,139,102,108,105,112,175,160,100,155,173,135,118,106,99,97,106,109,109,111,108,105,110,131,214,130,90,103,110,105,91,96,107,106,109,103,131,186,135,138,217,153,100,111,97,86,79,97,167,141,106,109,106,76,167,197,109,102,106,97,96,107,105,119,218,170,110,113,118,182,132,103),
(109,76,88,193,147,112,72,125,238,138,97,106,107,110,170,157,98,155,175,129,123,111,80,82,108,109,104,106,110,110,104,130,230,135,72,102,109,114,78,77,107,106,113,104,135,187,142,140,212,154,99,114,100,83,71,87,186,152,101,112,101,58,186,215,107,102,104,79,79,109,109,118,232,178,101,104,126,184,137,100),
(120,94,95,154,135,111,84,123,185,122,106,108,109,108,152,147,120,153,154,129,127,110,81,85,116,110,107,109,111,111,115,130,193,123,70,112,115,116,90,99,119,108,113,107,124,159,137,138,205,150,104,110,92,81,82,101,161,133,101,117,102,80,151,164,108,106,104,86,95,110,107,122,193,168,118,104,126,163,132,105),
(112,111,105,74,90,104,117,102,76,97,113,111,112,108,76,113,219,117,68,114,115,112,110,114,115,105,112,110,102,108,158,156,62,98,110,112,110,103,141,149,152,121,107,106,99,80,96,117,174,135,103,111,107,109,113,106,74,96,116,112,104,113,92,81,104,117,116,108,112,105,111,106,54,134,238,136,92,74,93,111),
(108,108,98,76,96,116,110,95,70,98,113,108,110,108,77,120,220,126,71,111,113,105,112,110,110,108,107,112,111,110,176,163,74,95,111,107,113,108,136,149,149,127,113,114,94,74,100,131,178,148,107,111,110,110,111,104,66,89,119,102,110,105,85,80,111,109,107,110,108,110,111,109,69,142,240,131,94,72,96,116),
(118,119,109,85,98,114,114,103,91,114,120,106,111,116,83,109,182,118,72,106,108,108,111,105,111,111,105,106,108,106,145,136,90,101,114,110,110,108,133,142,139,124,109,115,101,81,104,122,153,132,109,107,111,122,111,108,82,97,112,106,110,109,92,82,114,117,115,119,111,109,112,107,80,126,199,140,119,93,110,109),
(132,135,127,107,109,112,105,122,145,146,137,108,110,110,112,102,87,106,113,79,89,110,112,110,111,109,107,111,116,110,89,97,149,147,137,110,109,108,113,107,106,109,107,108,107,103,106,101,88,96,110,108,118,148,121,113,105,108,112,114,109,108,107,110,110,123,148,147,134,109,109,112,114,99,80,152,165,147,120,103),
(134,137,129,113,107,108,110,125,156,145,140,109,106,104,112,96,64,101,112,76,94,112,107,109,108,107,108,107,111,112,70,82,147,144,149,108,106,106,105,108,111,114,113,111,111,109,107,106,69,87,109,108,122,156,127,108,110,110,111,111,108,108,113,114,105,125,149,149,140,107,111,113,113,93,65,163,181,148,120,108),
(132,135,128,115,114,108,120,120,136,135,138,112,112,119,118,104,92,106,109,79,100,113,109,115,113,114,113,110,110,113,100,99,151,143,130,111,108,111,111,112,107,101,100,105,104,116,106,92,79,100,112,106,119,140,124,115,115,115,110,108,109,110,109,110,119,134,144,151,142,106,111,113,116,96,86,145,154,148,126,110),
(134,134,130,111,110,109,148,139,104,105,109,102,132,155,143,144,156,126,102,75,92,111,107,118,147,155,140,114,107,112,143,151,143,122,108,111,113,116,110,103,82,75,76,72,87,114,88,76,78,99,112,115,104,105,133,147,148,130,108,111,111,108,110,113,134,134,130,141,131,108,110,108,107,124,157,85,78,150,123,108),
(135,134,130,111,107,111,140,138,110,109,111,106,129,149,140,143,148,122,101,76,95,115,109,117,143,148,144,105,109,108,135,148,147,124,103,109,107,110,109,103,76,79,82,73,93,120,83,75,70,97,117,108,111,106,131,149,151,131,108,110,111,106,111,121,134,132,136,147,135,106,107,111,106,124,154,81,89,153,123,106),
(126,127,124,109,115,120,138,132,106,109,109,109,128,147,147,148,147,122,102,78,94,105,113,122,137,138,138,119,118,109,127,131,139,121,114,119,112,106,112,104,87,85,83,90,93,110,102,97,81,96,104,110,111,107,125,135,135,120,112,107,109,109,100,106,117,124,128,134,133,119,111,108,107,124,133,104,98,145,124,107),
(109,111,112,105,121,133,132,123,107,109,109,106,128,145,135,134,131,117,104,78,79,80,103,107,113,112,111,145,130,106,86,81,109,127,142,135,121,109,110,110,114,91,77,113,113,108,138,140,112,89,73,105,109,110,111,111,111,111,113,107,109,111,90,78,81,97,110,107,121,138,118,112,107,107,101,138,137,137,119,110),
(103,107,109,106,122,136,132,122,109,110,109,103,129,148,133,136,134,119,103,78,76,76,104,110,108,108,110,156,132,109,82,73,109,120,135,136,126,108,108,112,118,91,72,106,110,105,137,139,116,94,71,106,114,114,112,109,109,109,111,109,109,112,87,72,76,98,108,103,115,136,119,111,113,115,106,129,130,134,119,111),
(107,111,113,109,123,131,136,129,109,109,110,108,125,142,134,135,136,122,102,89,84,86,104,115,112,110,110,133,121,103,97,95,108,120,129,133,126,107,110,112,108,93,84,110,109,110,138,140,109,95,86,98,101,97,109,109,111,111,109,110,110,110,95,86,74,92,112,110,110,123,120,116,103,102,111,119,125,139,120,109),
(107,110,110,110,127,131,133,131,106,108,109,108,104,107,126,129,131,120,103,112,113,115,112,109,110,110,107,109,92,70,136,145,106,110,114,128,126,111,110,108,105,112,110,111,110,113,134,139,110,113,118,79,76,72,101,103,107,113,109,109,111,106,112,113,79,94,109,107,113,112,122,132,72,88,114,107,114,138,119,108),
(110,109,112,112,125,138,135,126,107,112,109,111,113,111,133,138,138,120,104,109,107,107,109,110,110,110,107,112,97,79,134,138,105,112,113,130,124,107,103,103,112,112,106,110,110,109,134,146,109,107,112,80,82,80,104,113,115,114,110,112,112,108,111,110,70,94,113,109,109,111,128,128,79,90,113,110,115,132,117,108),
(113,104,104,109,113,116,126,118,104,112,111,104,104,104,125,129,128,116,105,109,108,107,108,109,109,109,107,111,96,77,131,135,108,111,111,124,114,94,114,119,122,115,106,110,110,109,137,145,122,111,105,89,88,82,97,102,112,113,111,120,116,109,112,111,90,98,102,111,111,114,121,114,83,92,114,110,114,124,114,109),
(109,90,85,108,98,82,105,113,106,110,104,79,73,76,109,116,111,109,107,110,110,110,108,109,109,109,107,111,97,73,110,116,108,113,112,116,104,79,124,136,130,118,107,109,109,109,134,145,145,126,104,113,102,80,84,85,105,110,111,129,121,110,111,111,114,99,79,105,116,132,101,82,77,93,113,109,111,116,112,109),
(118,84,72,115,91,68,105,115,107,111,106,80,76,79,107,110,105,105,109,110,109,110,105,106,105,107,107,111,97,72,102,109,111,110,109,112,100,73,118,137,135,121,108,109,109,112,143,153,153,135,104,120,101,76,76,83,110,106,111,137,125,110,109,110,118,94,67,105,121,143,92,68,76,87,110,108,109,111,110,109),
(105,91,90,107,96,84,108,113,106,109,104,88,82,80,107,111,108,106,110,110,111,107,118,118,120,118,109,113,94,77,110,107,108,105,107,113,98,72,118,137,139,119,106,110,106,98,119,127,135,122,108,112,99,85,86,88,106,105,112,136,131,119,113,109,104,96,81,110,117,127,101,87,92,93,113,111,109,109,109,109),
(67,104,115,71,98,110,108,112,109,107,109,115,95,78,107,109,110,108,110,107,108,109,145,150,153,125,107,114,96,76,106,111,106,108,106,114,100,74,120,137,138,120,106,112,98,70,70,72,108,107,110,108,111,112,115,111,109,111,112,125,136,137,118,105,109,113,115,109,106,111,110,114,116,111,108,108,108,109,109,109),
(75,101,103,74,94,108,112,113,110,108,106,112,91,76,107,107,111,113,110,109,107,112,148,151,149,114,103,113,96,76,99,109,109,107,106,110,99,74,122,134,133,119,106,111,101,71,81,88,110,110,109,107,110,110,105,108,113,110,113,129,135,138,117,109,116,114,107,106,112,111,107,109,113,112,108,108,110,109,109,109),
(91,102,106,92,101,107,120,119,109,110,108,112,96,77,106,108,111,108,110,131,116,110,124,131,143,130,122,112,99,90,103,107,124,123,129,114,95,74,112,119,124,115,108,111,98,73,88,95,110,107,108,110,107,110,108,108,109,110,113,136,139,135,119,110,98,106,107,109,109,109,112,111,111,114,124,123,122,110,109,109),
(108,110,111,104,113,114,129,125,109,110,110,113,91,76,106,111,110,108,111,146,129,107,109,117,148,146,139,109,108,106,109,119,148,146,146,116,97,76,80,87,115,111,109,111,100,79,106,115,110,109,109,109,107,107,107,107,109,109,109,140,142,134,117,107,78,94,108,110,113,109,110,108,108,121,135,138,130,110,109,109),
(111,110,109,113,111,111,133,128,110,107,106,109,90,71,107,109,109,113,106,145,131,105,107,121,156,152,146,111,112,111,107,123,152,143,138,114,98,73,75,83,108,107,107,111,98,72,95,105,105,104,107,108,108,111,109,106,114,110,110,141,145,130,119,107,75,93,108,110,110,109,109,109,105,122,137,140,128,110,109,108),
(110,109,108,107,107,108,125,124,119,108,109,125,105,85,108,110,109,112,120,147,129,107,108,115,128,137,131,114,112,110,107,113,132,135,141,115,103,88,92,94,111,113,110,113,97,86,109,120,120,120,121,110,107,98,107,107,109,112,110,136,145,138,118,105,76,95,110,108,104,107,110,109,111,116,126,126,124,120,117,112),
(109,109,108,108,109,112,110,119,133,115,113,151,133,112,110,110,114,136,150,151,129,109,110,112,106,103,102,110,110,110,109,107,100,133,150,111,110,112,113,109,111,113,107,108,114,112,132,141,137,141,142,117,101,74,104,110,105,112,110,140,148,150,117,104,78,93,110,108,109,108,111,109,111,110,109,103,114,132,121,111),
(109,109,109,109,110,113,104,116,139,122,115,148,127,109,109,106,113,135,146,150,128,109,112,111,114,113,111,109,103,111,108,109,112,132,137,106,105,104,104,106,108,105,107,112,111,112,125,134,131,133,134,117,100,74,110,117,112,109,113,144,145,146,119,102,78,91,111,108,112,107,105,109,109,106,111,109,121,138,118,104),
(108,109,110,109,108,110,108,116,137,119,115,149,130,109,109,105,94,134,148,131,119,108,111,111,110,103,98,98,102,112,108,108,105,131,147,128,120,109,108,114,121,112,108,106,105,113,118,126,132,128,124,117,108,92,95,97,106,107,113,129,132,132,113,91,76,92,113,107,116,128,124,125,127,117,106,109,111,131,117,109),
(108,109,110,109,109,110,111,116,134,114,114,147,128,105,108,104,75,123,144,107,108,109,108,107,113,88,74,77,94,113,108,107,109,130,150,146,130,111,110,116,135,122,108,109,112,112,113,119,132,121,110,108,112,111,82,85,111,107,109,110,107,112,94,79,74,91,110,108,121,147,145,144,150,135,108,112,109,113,107,106),
(109,109,109,108,110,110,109,114,133,115,111,148,127,102,112,102,72,126,153,111,111,112,112,108,113,91,75,75,88,114,111,109,107,133,149,149,134,109,109,115,135,120,110,112,111,112,114,117,134,127,112,109,112,111,83,80,114,107,108,107,107,111,90,71,73,93,110,106,117,146,144,143,150,135,106,109,109,108,109,109),
(109,109,109,109,109,110,118,119,125,113,112,141,133,123,116,103,80,106,120,100,102,111,112,109,99,89,80,95,96,112,110,109,107,124,128,128,122,110,109,115,135,125,117,112,112,109,106,115,126,121,109,111,108,98,91,92,111,108,110,109,109,110,100,89,90,102,110,107,113,129,141,139,133,121,105,110,109,109,109,109),
(109,109,109,109,109,110,132,128,114,111,117,147,153,145,117,99,74,81,71,76,96,113,105,98,72,81,82,111,111,108,104,109,109,105,106,105,106,109,109,115,137,135,131,112,110,109,108,112,112,111,109,112,95,72,104,116,110,108,111,110,110,109,111,115,110,111,109,109,109,107,137,145,108,105,108,109,109,109,109,109),
(109,109,109,110,108,110,134,125,107,109,117,145,143,143,117,96,72,77,74,71,91,111,107,104,73,76,76,107,115,108,106,107,109,107,112,111,112,111,109,115,137,134,133,118,112,114,117,112,105,107,110,115,99,70,104,110,107,111,109,111,114,109,107,106,105,108,110,110,111,104,133,147,109,110,111,108,109,109,109,108),
(109,109,109,111,109,108,122,116,106,108,112,130,140,149,113,100,96,90,93,96,105,111,108,102,98,98,95,106,109,111,114,108,108,111,110,110,108,110,109,115,136,126,120,103,94,96,106,112,110,111,112,110,108,96,106,114,107,111,107,110,111,111,109,108,109,109,110,110,111,108,120,128,113,109,109,110,109,108,108,108),
(110,109,108,110,108,109,113,111,106,110,108,105,128,151,111,110,113,109,113,109,108,109,110,110,109,111,112,112,107,110,112,109,110,112,108,108,109,105,104,112,138,119,101,80,77,78,99,109,113,113,108,110,111,111,109,110,111,107,107,111,111,109,110,110,110,109,110,109,107,109,110,108,108,105,110,112,109,106,109,111),
(109,108,108,110,112,116,109,107,110,109,109,105,126,148,109,107,109,109,109,109,110,108,110,113,110,108,111,111,110,112,112,115,106,106,110,108,109,109,110,118,137,121,109,79,80,79,100,113,112,115,108,108,109,107,111,112,109,108,111,108,110,108,108,110,110,110,110,109,107,109,110,109,108,106,110,110,112,108,110,111),
(109,108,107,112,106,94,106,111,110,109,109,108,129,148,111,107,109,109,108,110,112,110,95,99,111,110,111,110,109,112,97,96,107,110,110,108,109,111,124,124,125,115,110,97,86,72,103,107,92,104,109,109,109,108,110,110,111,102,92,107,111,108,108,109,109,109,109,108,107,109,110,109,108,107,111,95,97,111,111,112),
(108,107,106,112,94,71,106,117,109,109,110,110,131,147,115,112,113,110,108,109,111,112,80,83,110,112,112,110,107,111,82,78,112,114,109,108,109,110,133,127,109,108,109,118,100,74,105,103,73,93,111,111,110,109,107,107,114,94,73,107,112,109,109,108,108,109,108,106,107,109,110,109,109,108,110,82,81,113,112,113),
(108,108,108,112,92,81,109,110,110,108,110,108,127,141,113,110,108,109,109,109,110,111,82,86,113,111,113,111,109,113,85,88,111,109,110,108,109,111,130,130,105,113,111,106,101,78,101,112,79,98,114,112,112,111,111,110,113,97,83,105,113,111,111,108,108,109,108,107,108,109,110,109,109,109,111,86,87,113,112,112),
(109,101,97,98,89,76,120,116,109,109,110,107,116,132,102,97,104,108,110,108,108,112,76,80,111,112,114,109,103,99,76,86,125,112,109,109,109,108,120,117,93,103,108,106,108,93,107,108,72,92,113,114,114,107,98,97,99,85,78,115,118,108,109,108,108,109,107,103,104,111,109,108,107,109,111,80,78,112,116,118),
(116,85,76,78,77,82,130,123,108,109,109,110,109,106,79,85,109,108,111,109,107,110,82,86,113,124,128,115,95,76,77,94,136,115,108,109,109,106,112,102,75,93,109,109,113,112,110,103,74,97,114,130,123,113,85,75,78,81,80,123,126,110,110,108,108,111,110,79,82,112,109,103,111,108,105,87,81,115,126,135),
(111,82,74,80,78,76,130,130,107,109,109,109,108,107,80,88,116,115,113,111,106,113,77,80,109,127,134,122,94,75,74,88,140,120,107,109,109,109,111,100,79,99,117,115,111,110,108,107,69,91,113,133,131,117,82,75,78,73,78,126,125,112,110,108,109,109,110,83,87,114,117,114,113,107,109,83,78,110,122,133),
(107,100,96,96,93,97,119,116,109,109,109,110,109,106,83,84,91,94,95,111,108,109,94,99,108,118,118,111,103,94,92,100,123,113,109,109,109,106,108,101,74,85,94,91,100,110,107,108,93,104,109,122,115,109,97,96,95,94,96,121,119,109,109,108,109,109,111,81,81,98,93,94,111,110,110,98,94,111,118,121),
(112,112,112,112,111,115,107,105,110,109,109,108,108,110,84,76,73,75,78,111,111,107,110,114,108,109,106,103,111,112,113,112,105,107,110,109,109,111,110,103,78,75,73,71,87,116,108,107,113,113,107,111,103,104,113,113,109,117,113,108,112,108,111,108,108,110,110,86,80,80,70,79,107,108,109,112,109,109,112,109),
(108,106,106,113,110,109,110,114,111,110,109,108,110,105,80,79,81,80,78,112,108,107,109,110,106,111,110,111,107,111,107,109,111,114,110,110,109,111,112,100,75,79,82,76,86,113,106,107,111,108,107,111,110,109,108,111,110,103,107,112,107,110,114,111,111,110,108,84,78,80,77,82,108,108,106,106,108,111,110,109),
(108,109,112,114,108,112,109,113,113,95,91,109,111,109,99,91,74,93,95,108,119,127,112,110,110,100,94,117,117,112,110,110,110,114,110,90,96,110,110,107,98,85,78,95,98,112,123,124,109,110,109,93,100,120,111,107,113,114,106,105,111,112,98,98,111,110,111,103,94,77,94,97,109,116,127,115,109,110,94,84),
(108,109,110,105,108,112,107,111,112,85,79,108,108,111,114,101,76,103,114,108,127,146,114,105,113,87,80,107,108,105,110,111,107,113,107,78,88,111,108,112,113,91,80,111,112,109,137,140,107,109,110,79,89,112,111,106,105,109,107,110,111,113,83,73,110,109,107,112,107,78,104,120,108,124,152,117,108,114,92,75),
(108,109,109,115,115,110,104,101,108,87,82,106,109,108,109,101,71,93,106,100,125,157,115,107,113,87,77,105,108,117,113,108,101,104,104,81,89,109,109,107,110,91,72,100,106,100,142,147,108,109,110,78,87,110,109,116,117,108,109,105,100,106,84,76,112,110,107,109,101,71,93,105,102,126,153,121,106,110,93,81),
(108,110,107,92,106,111,127,127,133,100,93,109,109,108,108,109,95,119,129,127,126,120,109,108,110,91,83,109,100,95,109,115,128,129,128,92,99,110,108,107,110,105,97,127,127,128,125,117,108,108,109,83,91,110,110,110,95,97,112,123,126,129,105,94,111,111,107,109,107,93,116,131,135,127,123,110,109,109,91,79),
(109,109,105,74,97,108,143,148,152,124,111,111,107,111,115,110,106,136,152,151,128,106,111,107,111,91,82,111,99,76,102,115,150,148,148,115,112,110,107,114,113,109,109,147,150,150,116,109,110,108,109,82,90,112,111,100,76,91,112,142,150,154,127,114,107,109,110,108,111,113,138,148,150,128,108,106,109,108,90,79),
(108,111,106,77,93,110,141,142,147,123,106,112,110,109,110,107,109,137,150,145,128,110,109,106,112,87,79,112,98,77,101,117,146,141,146,113,108,112,109,110,109,107,113,145,147,144,120,110,107,108,109,78,87,113,114,107,80,92,111,140,145,144,118,107,106,112,112,110,106,108,138,145,144,131,104,109,108,110,87,76),
(108,104,94,77,91,113,126,131,143,118,110,112,107,107,110,110,108,123,129,145,129,108,108,113,133,96,80,114,98,74,103,116,128,135,140,111,113,110,107,108,110,110,110,127,131,147,118,109,107,120,129,82,89,113,99,95,81,97,111,122,136,146,122,108,110,110,111,110,110,104,120,131,146,131,110,108,111,134,97,76),
(110,83,73,77,101,111,105,122,149,114,104,107,111,112,107,108,105,105,112,143,129,107,109,119,152,104,77,113,96,76,109,114,105,133,145,105,107,107,112,110,107,108,104,106,119,146,118,108,108,130,148,85,89,114,81,76,78,98,109,103,112,148,122,108,109,108,106,105,112,112,106,110,147,131,105,107,116,153,102,75),
(115,82,74,67,89,110,100,125,154,119,104,107,111,117,116,116,114,115,114,143,129,107,108,116,151,100,76,112,94,73,99,105,102,138,148,110,106,108,113,117,115,115,114,113,121,146,118,108,107,127,147,82,88,116,85,74,73,95,114,109,120,155,127,106,112,114,113,112,113,116,112,113,143,132,110,108,115,150,102,77),
(112,99,97,95,103,110,110,116,126,118,106,114,101,91,93,91,92,91,95,146,130,106,110,121,153,102,78,112,106,99,108,109,111,120,126,113,106,114,95,92,92,90,94,88,108,149,118,107,110,131,149,83,87,116,107,99,97,101,113,111,111,124,115,107,110,96,93,92,88,90,92,101,144,131,108,106,117,154,107,75),
(112,115,112,111,110,109,113,108,103,104,108,115,89,70,77,76,78,69,79,145,129,107,105,114,150,102,80,109,111,111,110,111,111,107,101,106,109,114,75,72,78,78,80,66,101,151,118,107,104,125,148,85,87,112,110,109,113,110,109,108,107,104,107,109,112,88,75,78,74,74,74,84,145,129,106,107,115,154,100,69),
(107,107,105,107,108,107,107,111,112,112,112,112,98,82,80,77,78,77,88,144,129,107,109,119,149,104,79,105,109,109,111,108,107,112,112,112,111,111,88,80,78,77,81,78,102,149,118,108,110,128,147,86,92,110,111,112,110,111,108,108,112,113,113,110,112,95,80,77,79,78,74,83,145,128,106,108,118,152,102,73),
(110,109,111,112,112,110,109,104,92,111,110,109,104,98,98,97,97,96,105,146,130,108,109,114,128,109,97,111,110,106,110,108,110,98,96,113,108,110,100,96,97,98,99,95,110,145,120,107,110,117,128,100,103,113,110,108,108,106,104,112,104,88,104,111,109,106,96,114,121,129,110,97,140,127,107,108,113,130,110,95),
(106,106,107,111,112,108,110,100,71,105,109,111,107,110,115,113,113,109,112,135,128,109,106,105,104,111,111,112,109,106,110,106,112,88,77,111,108,111,106,111,113,112,111,104,124,146,119,107,106,105,106,113,112,116,110,105,111,113,109,114,103,69,98,112,108,112,108,142,149,150,126,118,137,129,109,108,106,109,117,116),
(109,114,113,111,110,107,112,102,74,97,114,114,110,111,111,110,109,107,115,133,120,109,111,111,107,111,112,112,109,111,110,106,114,92,77,105,115,113,110,108,102,100,104,105,119,134,115,109,112,110,107,111,112,112,116,114,114,112,110,110,104,75,98,111,108,104,106,138,146,155,121,112,133,124,109,109,108,109,110,108),
(106,93,81,89,103,110,116,104,98,102,111,111,110,107,109,109,110,108,110,121,113,108,113,112,110,107,108,111,106,85,100,113,114,100,98,104,112,110,108,116,136,135,132,112,107,117,110,110,113,111,109,106,109,107,92,91,87,92,110,111,104,101,110,109,108,123,134,149,142,121,112,108,117,111,108,109,110,109,104,109));

CONSTANT BASE_B: my_background :=
((35,32,33,31,34,35,34,41,36,29,35,37,38,26,26,31,29,32,45,21,20,23,29,37,34,32,31,39,35,27,26,31,26,26,27,41,34,33,30,32,39,34,29,34,36,32,27,32,39,38,25,21,21,35,36,35,32,31,18,28,27,35,23,38,24,29,29,28,35,35,35,31,25,34,40,39,25,31,33,31),
(33,24,24,31,20,19,27,27,18,23,32,21,21,23,29,28,30,30,18,26,35,27,23,22,17,26,30,24,30,25,26,22,19,32,35,22,21,31,23,24,24,25,28,32,28,19,33,39,17,23,18,36,32,31,31,28,25,19,22,40,37,23,23,30,18,32,33,23,31,32,26,21,38,31,19,21,20,26,29,32),
(29,27,22,20,30,24,81,67,20,27,31,27,23,33,87,70,34,22,27,89,63,30,25,26,26,66,91,29,25,29,20,29,21,69,91,24,23,33,27,27,19,65,92,36,24,23,82,81,18,22,32,97,80,22,21,19,24,23,38,80,70,15,21,30,26,29,26,77,79,29,21,36,94,58,19,27,26,28,29,30),
(20,24,20,3,26,34,93,77,21,29,26,28,25,32,103,78,12,1,20,106,57,9,14,24,19,69,100,39,30,23,9,24,23,82,93,17,24,29,25,26,17,72,100,28,7,15,83,85,23,19,25,94,77,19,25,10,13,24,37,96,65,21,20,26,26,25,21,89,86,16,6,31,96,63,18,25,20,28,26,25),
(39,30,21,33,27,24,77,62,10,41,40,19,20,25,74,69,27,37,47,76,52,20,30,30,15,68,76,25,17,24,40,37,14,55,77,43,35,39,24,21,17,56,79,34,23,40,67,71,27,18,20,76,62,34,38,22,39,34,16,68,67,31,37,34,16,34,36,70,65,24,29,47,73,57,23,22,27,45,31,19),
(86,36,16,93,46,5,40,27,7,72,77,15,19,18,28,33,29,82,97,20,25,33,22,24,23,24,23,25,17,22,76,70,12,29,44,74,83,85,29,18,30,30,29,28,53,87,46,26,25,22,19,28,48,86,47,36,93,52,6,28,36,48,80,86,20,33,47,31,31,30,64,71,32,33,26,12,37,90,51,19),
(100,47,25,110,62,18,21,20,12,81,87,22,22,15,14,16,22,72,82,7,27,20,14,25,32,13,16,22,22,38,87,87,24,19,17,81,98,105,36,11,23,20,11,32,61,99,40,15,29,27,25,15,50,109,51,34,101,54,7,18,31,55,91,84,15,38,59,22,20,17,71,95,23,20,29,15,37,102,57,20),
(91,53,33,90,53,25,21,20,20,70,78,21,9,13,29,35,16,60,82,28,35,28,22,22,39,30,31,24,19,38,69,71,27,20,23,95,99,83,37,19,25,26,31,25,43,82,40,22,28,24,25,22,46,94,44,31,80,56,22,24,32,57,90,91,22,38,64,38,33,12,78,106,16,14,28,21,38,85,52,24),
(67,65,51,24,16,17,21,14,16,18,27,27,36,36,46,41,36,42,50,47,36,36,24,34,96,43,19,26,21,23,23,16,8,30,43,45,27,21,20,32,27,34,45,20,18,22,23,24,29,22,22,22,18,20,22,33,34,23,17,19,41,91,49,57,25,48,89,49,32,27,38,36,22,19,27,20,18,30,22,17),
(57,53,42,13,18,31,27,23,27,13,19,21,16,15,49,45,31,43,60,60,45,27,19,31,106,59,29,26,16,29,23,27,22,29,24,63,39,22,23,20,16,44,68,25,15,24,19,22,30,22,23,28,32,26,17,32,26,30,26,15,39,85,59,47,29,53,85,59,45,31,42,46,24,25,39,26,23,37,35,27),
(52,63,63,30,34,38,19,23,47,20,24,46,38,29,50,49,11,44,58,58,55,33,32,47,93,51,23,25,28,30,24,36,46,25,17,65,41,31,44,28,36,42,42,38,29,20,16,20,24,19,29,38,36,31,19,24,29,28,30,14,36,78,59,42,34,54,78,63,48,10,55,68,18,31,39,18,22,39,35,43),
(74,81,86,85,74,41,24,23,42,31,38,54,46,41,63,54,17,89,117,115,92,38,83,73,30,43,61,13,36,63,53,45,46,28,24,59,52,22,62,38,45,48,43,25,28,20,16,15,29,22,25,48,32,18,24,25,34,47,52,22,30,94,50,32,52,72,72,94,72,22,71,99,27,34,48,32,45,95,49,40),
(80,74,74,97,81,62,32,29,57,32,29,56,68,65,62,41,25,93,118,113,97,45,106,72,27,40,48,20,39,65,56,63,63,33,26,55,47,16,54,64,49,60,58,27,23,20,28,25,32,16,25,38,48,35,16,32,70,72,66,22,38,87,41,33,49,64,77,82,73,25,78,115,38,46,59,32,34,109,67,52),
(66,60,75,105,55,46,31,30,60,42,32,41,56,57,65,48,27,86,110,109,90,45,93,74,41,51,54,19,37,56,56,47,57,41,32,54,41,26,37,48,50,57,53,44,33,17,41,48,26,17,35,44,47,30,18,30,61,50,51,32,37,74,31,34,58,77,77,60,57,25,93,114,28,43,51,24,49,83,62,55),
(149,63,16,50,73,80,17,36,93,62,58,78,67,68,99,86,45,66,86,110,87,72,30,33,39,67,81,46,68,86,81,74,83,49,6,46,73,58,42,27,69,85,71,45,34,21,38,29,23,51,61,81,58,10,10,27,72,84,92,63,49,5,55,58,79,59,73,42,36,67,54,67,25,45,88,62,53,24,52,79),
(143,54,12,55,80,79,34,52,74,58,57,71,78,71,94,83,42,68,92,107,89,67,34,40,67,67,81,54,59,74,73,79,83,48,28,59,62,48,19,43,66,84,77,59,54,16,52,56,20,42,63,69,67,29,17,31,82,81,68,65,41,18,47,67,69,71,62,19,30,55,81,95,27,41,86,61,30,9,48,76),
(131,52,28,45,66,75,40,51,77,70,59,68,66,70,78,70,63,55,67,121,95,65,43,45,51,66,66,68,75,80,72,77,70,45,50,62,61,41,37,52,74,76,80,56,42,16,77,74,27,55,57,63,61,48,26,45,68,78,69,65,56,29,43,40,70,69,70,46,45,53,70,88,51,53,73,66,42,20,57,80),
(87,57,47,38,59,76,43,32,33,72,75,74,69,69,37,39,84,46,44,129,106,84,53,50,81,73,74,83,84,78,82,82,25,41,45,73,88,90,48,52,70,71,80,98,66,11,105,114,22,57,79,81,69,44,55,43,40,56,77,82,72,49,28,29,79,74,66,56,54,79,77,80,84,79,64,79,72,27,58,75),
(67,68,61,20,43,83,64,46,1,54,80,77,73,70,39,43,81,48,34,149,112,81,64,64,82,70,75,74,78,82,87,64,2,51,65,71,79,89,71,62,66,72,80,85,66,26,113,115,5,44,78,76,68,58,71,44,18,48,85,73,78,67,26,24,72,72,72,62,60,84,78,73,95,96,74,80,64,22,52,76),
(78,63,47,33,63,80,56,54,27,66,85,77,75,76,41,45,78,54,43,132,98,70,60,65,83,71,76,74,80,80,65,58,26,56,59,81,79,74,63,65,77,76,76,71,61,40,105,106,17,49,81,73,63,54,47,47,39,60,78,79,72,44,43,49,69,67,76,48,57,83,74,81,94,91,74,80,63,32,57,80),
(86,80,79,40,71,75,76,64,49,76,80,75,74,81,53,41,24,42,64,64,85,83,82,81,81,74,73,74,85,82,45,37,54,58,81,90,77,74,102,107,113,90,73,82,69,25,75,79,8,54,79,73,83,80,85,93,51,64,77,82,74,85,55,39,69,76,79,82,82,70,81,72,26,64,104,82,82,54,61,69),
(72,74,82,45,70,73,70,74,57,71,87,78,75,71,54,50,15,41,61,88,82,78,82,77,77,76,75,76,85,73,34,25,55,72,76,76,80,82,103,112,117,97,81,85,77,59,73,62,32,60,82,75,78,76,76,78,50,65,80,79,81,89,66,62,88,90,75,80,76,75,78,74,65,65,96,70,70,54,69,79),
(95,95,96,52,70,74,78,77,64,83,90,74,78,77,65,59,37,51,63,76,78,79,81,72,78,78,74,70,77,74,48,38,70,75,81,76,77,78,101,106,106,91,76,80,78,62,79,66,47,67,87,73,77,88,71,72,54,71,76,83,83,81,73,64,79,84,82,84,76,75,78,72,64,70,96,58,72,68,78,77),
(131,128,118,77,81,76,68,85,109,112,102,75,76,75,83,68,48,63,89,51,59,81,82,76,78,76,74,76,84,88,50,61,119,113,107,77,76,76,79,73,72,75,73,71,76,73,82,71,35,66,89,73,85,114,87,79,72,82,79,87,81,81,79,71,68,85,110,112,100,75,75,81,82,70,49,31,51,120,88,69),
(139,138,123,84,76,74,73,86,118,111,105,75,72,69,79,69,60,69,78,52,63,84,77,75,74,72,75,74,77,89,56,70,111,109,117,74,74,72,71,77,80,83,82,78,79,74,79,89,46,67,82,74,89,122,93,73,74,83,82,82,81,79,80,78,76,95,114,114,106,73,77,82,73,76,50,36,30,111,87,75),
(125,133,121,83,79,74,83,87,104,101,105,79,78,83,83,71,55,70,68,61,68,85,79,79,79,78,79,78,76,80,76,76,111,117,96,78,74,74,78,85,80,74,73,79,75,77,73,75,58,67,72,73,86,105,88,79,80,85,84,81,83,79,72,81,99,109,115,117,107,73,77,77,76,73,62,45,55,114,90,77),
(132,136,125,82,76,76,111,107,75,76,80,73,100,118,108,112,112,87,68,53,63,81,74,84,113,121,106,81,73,77,104,121,113,86,70,77,83,84,78,74,55,50,51,47,59,82,57,56,55,67,77,81,72,72,98,112,113,97,78,80,83,79,76,83,122,129,116,109,92,68,74,84,74,92,114,56,61,114,85,77),
(135,132,122,84,78,81,107,107,79,83,84,79,98,115,100,109,112,87,76,51,71,86,75,83,109,115,112,72,77,75,98,116,120,92,70,73,74,81,80,72,47,54,59,46,64,92,56,52,47,74,91,73,78,73,97,115,117,97,73,76,81,78,80,92,125,135,129,118,96,73,74,88,77,89,110,61,66,116,91,76),
(115,115,107,82,89,99,118,108,75,83,82,81,95,114,114,120,117,94,78,57,75,80,82,88,103,105,106,86,86,79,103,98,104,110,98,92,80,77,83,73,59,58,59,62,64,80,74,72,55,70,78,76,76,72,91,102,102,87,78,74,80,80,70,81,102,112,115,108,100,112,86,68,74,90,104,84,84,129,99,73),
(92,92,86,75,101,123,125,106,76,83,82,80,94,114,123,135,127,97,80,57,61,57,74,73,79,78,79,112,97,78,66,54,78,115,140,130,106,81,80,79,85,64,51,85,82,76,109,111,80,62,47,73,74,75,78,78,79,77,79,73,79,82,61,55,60,75,87,81,94,143,98,71,76,73,85,132,137,131,101,74),
(75,75,71,72,109,140,138,113,79,83,82,78,95,119,127,142,136,102,75,55,57,51,74,76,73,74,77,123,100,80,59,49,78,103,132,136,116,82,79,81,88,64,46,77,77,71,106,103,79,66,45,78,84,85,81,78,79,76,77,75,80,83,58,49,53,69,75,77,95,139,99,82,86,82,84,121,129,126,103,79),
(71,71,69,73,111,138,142,119,78,82,82,81,89,115,120,129,126,101,69,63,62,59,73,82,79,77,78,100,90,75,69,67,77,99,116,129,113,77,78,78,78,64,55,79,77,77,105,101,72,67,59,74,77,71,81,79,80,76,76,78,78,80,65,60,51,62,75,81,89,110,101,105,81,72,80,95,111,131,104,78),
(74,76,76,73,111,131,136,118,78,82,81,78,66,79,115,128,123,98,66,86,85,86,83,81,81,81,78,80,65,46,106,112,76,78,89,130,117,79,76,72,74,78,76,82,82,83,101,107,79,84,89,56,53,44,71,74,72,76,80,80,74,73,81,86,54,69,77,72,79,77,112,135,53,59,86,77,94,138,100,73),
(78,77,81,75,104,138,149,121,84,85,81,82,79,82,127,142,139,100,68,82,79,78,80,81,81,80,78,82,69,54,105,103,70,76,86,124,111,82,80,79,83,84,79,81,81,78,101,113,76,77,83,56,58,53,75,84,82,82,81,83,81,75,80,82,45,68,82,75,78,85,117,124,60,61,84,80,93,125,95,76),
(81,76,78,73,88,107,120,94,74,86,82,76,73,76,109,115,115,94,72,80,80,78,79,80,80,80,78,82,68,52,102,98,70,72,81,108,95,70,95,103,99,92,82,81,81,79,104,112,89,79,75,62,63,56,69,73,82,84,80,94,92,76,80,82,63,72,72,78,81,97,111,103,63,63,82,80,88,109,87,79),
(80,65,63,74,74,63,78,75,73,85,75,51,46,49,79,78,80,85,77,79,81,81,79,80,80,80,79,82,69,49,80,81,74,79,81,89,78,55,107,128,120,99,79,80,80,79,101,113,112,93,73,86,77,56,57,56,78,78,80,113,105,77,79,81,86,71,51,73,91,124,90,61,57,65,80,80,81,92,80,82),
(88,60,53,84,66,48,78,85,80,84,77,52,51,52,75,69,72,81,79,79,80,81,76,76,76,78,78,82,69,47,72,76,81,80,79,79,71,53,108,138,136,102,74,80,81,82,110,120,119,101,72,92,75,52,51,54,84,72,79,128,112,76,76,79,88,67,39,73,99,143,79,41,56,59,76,79,76,83,75,83),
(76,64,64,74,69,66,82,85,80,80,75,58,57,54,79,81,75,72,76,76,78,74,85,83,85,84,77,80,64,53,82,75,76,72,75,83,71,49,112,143,143,102,70,80,81,74,89,95,104,93,78,83,70,56,56,61,83,76,79,131,121,98,80,77,70,67,50,77,93,117,83,58,66,67,87,82,79,80,80,80),
(41,76,85,42,70,84,76,80,80,78,80,85,70,52,79,80,76,74,76,73,75,76,112,115,118,91,74,80,66,52,78,78,73,75,74,84,73,52,114,140,141,103,73,82,73,47,44,44,78,78,81,79,82,83,88,86,85,78,82,125,138,135,98,73,76,83,85,79,73,78,77,82,88,80,75,74,76,80,80,80),
(51,71,70,49,62,74,78,82,80,79,77,83,67,51,79,78,78,79,76,76,74,79,115,116,114,80,70,79,65,50,68,75,77,74,74,81,72,52,113,130,128,101,77,81,76,48,59,63,82,81,80,79,83,82,78,81,84,75,84,125,133,142,98,78,87,85,77,77,77,71,74,80,81,80,72,75,78,79,80,80),
(65,70,74,67,68,73,95,93,78,81,79,83,72,52,78,79,77,74,76,97,83,77,91,96,108,96,89,78,68,64,71,72,92,90,97,85,68,50,97,105,108,93,80,81,72,50,64,69,82,78,78,82,81,84,81,79,77,76,83,117,121,134,92,80,72,76,78,80,78,75,85,85,77,89,101,104,98,80,80,80),
(76,78,81,76,78,86,119,106,79,81,81,84,69,52,79,81,77,74,77,112,96,74,76,82,113,112,106,76,76,81,76,82,116,113,113,87,70,48,56,63,89,84,79,80,75,55,77,84,78,81,79,82,82,81,77,77,78,80,76,105,119,137,91,78,54,63,79,81,84,75,78,80,74,105,133,137,115,81,80,80),
(81,80,80,84,80,84,132,120,80,78,77,81,62,45,80,77,73,81,73,111,98,72,74,87,122,119,115,80,82,83,77,90,120,110,105,82,68,47,53,55,77,75,80,82,68,45,69,77,85,72,77,79,80,85,81,74,79,76,74,99,122,140,94,74,52,66,79,81,79,74,75,77,70,103,134,147,121,78,79,79),
(81,80,79,78,78,81,112,115,100,80,77,94,75,57,80,78,73,81,88,113,96,74,75,81,94,104,99,82,82,81,79,82,99,102,107,81,72,61,69,63,72,74,80,85,65,54,84,98,98,91,92,76,77,71,80,75,73,77,74,97,118,129,91,72,53,69,81,80,73,74,77,79,77,90,110,111,106,98,92,82),
(80,80,79,79,80,84,78,100,131,89,74,115,103,83,82,79,81,105,117,117,96,76,77,78,72,69,68,75,78,82,80,76,67,100,116,78,79,81,82,75,72,77,77,79,84,81,117,136,119,134,134,84,69,45,75,80,72,77,75,105,114,110,89,75,55,67,81,80,78,75,78,80,79,79,84,64,88,127,104,78),
(80,80,80,80,81,86,64,93,146,97,74,112,95,80,79,77,83,105,113,116,95,76,79,77,80,80,79,76,73,83,79,78,78,99,103,73,75,71,71,75,81,79,79,83,82,86,126,145,133,145,144,90,66,45,81,88,81,74,78,113,110,99,90,76,56,64,82,79,81,74,72,78,77,70,86,71,100,136,101,71),
(79,80,81,80,78,83,74,94,141,95,75,115,96,78,79,76,66,105,116,96,86,75,78,77,75,71,71,72,75,82,79,76,71,98,113,95,90,79,76,89,104,92,77,76,76,88,102,119,130,120,112,88,76,64,66,69,77,71,79,99,100,103,84,67,55,65,83,78,86,94,91,91,91,82,76,77,88,117,96,77),
(79,80,81,80,79,83,78,96,137,92,77,114,94,72,75,76,48,93,111,74,78,77,74,75,78,56,49,49,66,84,79,77,78,98,117,113,98,80,77,91,130,102,71,80,84,82,76,89,124,101,74,72,80,83,55,57,83,74,77,80,75,89,67,57,53,65,80,79,90,114,112,109,115,101,74,82,81,85,79,74),
(80,80,80,79,81,81,72,94,130,94,75,113,92,67,76,75,46,96,124,82,85,81,76,78,82,61,50,46,59,85,82,81,78,104,118,115,100,75,74,87,138,99,73,84,80,79,76,86,129,117,77,73,80,82,58,54,84,79,80,77,71,79,65,48,50,69,81,77,86,113,111,110,118,101,78,83,82,76,76,76),
(80,80,80,80,80,79,93,105,107,90,77,107,98,88,81,77,54,78,92,72,73,80,80,79,74,65,51,67,68,83,81,80,78,95,96,95,89,76,75,87,129,110,94,81,77,76,71,86,108,96,76,81,82,72,65,64,81,79,81,80,76,80,73,65,66,77,80,79,82,96,108,106,100,88,76,83,82,79,78,78),
(80,80,80,80,79,82,127,128,90,84,83,112,118,110,82,74,50,53,43,48,65,82,75,69,49,59,52,84,83,79,75,80,80,77,74,72,72,75,75,87,139,135,125,82,75,77,74,80,82,78,76,85,72,48,78,86,79,79,82,81,77,78,83,88,82,83,80,81,78,74,104,112,75,72,79,83,82,80,79,79),
(80,80,80,81,79,84,128,122,78,78,83,110,108,107,83,71,48,49,46,43,61,80,76,78,48,51,48,78,85,79,77,78,80,78,80,78,78,77,75,87,142,134,126,93,78,85,82,76,68,76,79,85,73,47,77,79,74,81,80,81,83,79,77,76,75,78,81,81,80,71,100,114,76,77,82,82,82,81,81,81),
(80,80,80,81,79,80,98,93,72,76,79,96,105,114,80,75,72,61,64,68,76,79,76,76,69,69,68,75,78,82,84,79,78,82,78,77,75,77,75,87,135,112,98,80,64,70,70,74,72,82,81,77,80,72,79,82,74,82,78,80,82,79,77,78,79,80,81,81,80,75,87,96,81,77,80,81,81,82,81,81),
(81,80,78,75,78,81,83,78,75,81,80,72,93,118,82,83,86,80,84,80,80,78,76,76,77,80,83,83,75,75,83,82,81,79,78,79,78,74,72,86,135,103,75,53,54,58,68,78,84,81,78,81,83,82,80,81,82,80,82,80,77,76,77,81,81,81,81,80,78,80,81,80,79,76,82,74,80,81,76,72),
(80,80,78,76,83,89,81,75,79,81,81,72,92,115,81,81,82,80,80,80,80,77,79,81,78,76,79,79,76,79,83,88,78,74,80,80,80,75,80,92,129,102,81,51,55,57,69,82,84,85,79,78,79,77,82,83,80,81,86,77,78,76,77,81,81,81,81,80,78,80,81,80,79,77,82,74,82,80,77,75),
(80,79,77,81,77,67,78,81,80,80,81,75,95,115,82,80,82,81,79,80,79,79,66,70,79,77,78,76,76,82,69,70,81,80,80,80,80,74,101,102,108,92,80,69,60,48,73,76,65,77,80,77,77,76,80,81,82,76,68,78,79,77,78,80,80,80,80,79,78,80,81,80,80,78,82,65,68,81,80,80),
(79,78,77,84,66,44,80,88,79,80,81,78,97,114,86,86,86,81,79,80,76,81,55,57,79,79,81,78,76,83,54,52,86,86,80,80,80,72,116,111,83,81,76,90,74,47,75,71,48,69,82,80,80,79,78,79,84,67,49,78,82,79,79,79,79,80,79,77,78,80,81,80,80,79,81,56,52,82,83,85),
(79,79,79,85,64,55,84,82,81,79,82,75,92,108,84,83,81,80,81,79,74,81,58,61,83,77,83,81,80,86,57,63,86,82,81,79,81,72,120,120,73,81,77,78,75,50,71,79,54,75,85,81,83,83,83,81,83,72,61,75,84,83,82,79,79,80,78,77,79,80,82,81,80,80,82,63,57,80,83,86),
(76,75,75,72,62,51,97,90,80,80,81,78,89,103,72,68,74,76,80,79,74,83,54,61,78,95,96,78,73,73,49,61,102,85,80,80,80,77,103,101,69,71,70,75,77,62,76,79,50,70,82,100,92,76,69,68,70,59,55,102,98,71,80,80,79,80,79,78,76,78,74,75,77,81,81,59,48,76,96,106),
(86,61,55,53,51,60,126,115,82,80,80,82,84,78,52,57,76,78,81,80,75,81,58,67,83,117,125,94,70,52,51,76,134,102,79,80,80,76,88,79,53,63,74,79,83,80,79,76,51,75,86,129,115,90,59,48,52,52,57,118,112,73,80,80,79,82,82,53,54,79,74,71,81,78,75,64,51,88,119,136),
(87,58,50,55,53,52,132,129,78,80,80,80,82,78,56,63,83,86,84,80,75,85,52,56,82,122,130,101,69,50,48,70,147,109,76,81,80,77,82,75,54,72,87,87,82,77,78,80,44,66,89,133,121,93,57,49,53,41,53,119,114,79,79,79,80,79,80,57,61,84,85,84,84,75,78,57,48,85,113,132),
(83,75,69,68,66,67,101,97,74,81,80,81,84,78,59,61,64,68,66,79,79,82,66,72,79,102,97,78,72,67,64,72,108,87,76,81,80,77,76,73,52,61,69,66,70,77,77,82,64,76,82,108,89,75,69,70,69,61,67,107,102,77,78,79,80,78,79,55,57,71,64,66,82,76,77,70,64,77,93,100),
(82,82,82,78,77,82,72,71,81,80,80,80,82,82,57,53,53,53,50,78,84,79,81,85,73,80,75,71,81,78,80,78,69,75,81,79,81,86,80,77,59,52,50,49,58,82,80,83,85,83,71,84,70,74,84,84,80,86,81,85,84,73,80,78,80,79,76,62,58,54,43,52,77,72,75,80,80,75,82,77),
(77,75,75,78,76,74,73,79,82,81,81,78,83,77,51,55,64,57,50,81,78,76,77,80,74,81,82,83,78,76,72,75,73,81,81,82,79,84,83,72,50,57,61,52,57,82,75,78,80,78,75,83,81,79,77,78,76,71,75,84,77,79,87,85,80,76,75,57,53,56,50,53,78,75,72,73,77,76,79,79),
(79,81,82,81,76,77,75,78,79,69,64,79,82,80,70,65,55,67,66,78,86,94,78,79,85,73,68,88,84,79,77,75,76,78,78,65,68,80,82,77,69,62,58,67,69,81,90,90,76,81,84,68,72,85,78,76,79,83,76,76,82,85,74,74,79,74,80,74,66,52,67,66,79,86,95,82,76,74,62,59),
(79,80,80,73,76,80,73,76,81,63,57,80,79,82,84,74,53,76,85,76,94,114,81,75,87,60,53,79,78,72,78,78,73,78,78,57,63,82,79,83,84,66,56,82,82,77,104,107,75,80,83,53,61,78,79,75,74,80,77,79,79,84,57,47,79,77,78,84,79,52,76,88,76,92,119,84,75,83,66,53),
(79,80,80,82,84,79,71,67,77,65,60,78,80,79,79,73,43,64,75,67,92,124,82,76,87,60,50,77,79,84,82,77,68,70,77,60,65,80,80,78,81,63,45,71,74,67,109,114,75,80,84,51,58,77,75,85,89,81,79,73,67,76,56,49,82,82,81,80,71,45,64,71,69,93,120,88,73,81,68,60),
(79,81,78,60,76,83,94,93,102,75,67,80,80,79,79,78,63,89,97,94,93,87,76,77,85,64,55,81,71,61,79,86,95,96,98,67,72,81,80,79,79,74,66,97,94,94,92,84,75,79,83,56,62,77,76,80,69,72,82,89,93,97,76,63,82,85,83,80,75,66,86,97,101,93,89,77,76,80,65,55),
(80,79,75,44,66,79,110,115,119,95,82,80,77,81,85,79,74,104,118,115,95,73,79,77,83,63,54,83,72,46,74,85,116,115,116,87,82,79,77,83,84,77,78,115,115,115,83,76,78,79,81,55,61,81,78,70,51,66,82,108,116,121,96,83,79,84,85,78,80,87,109,114,114,94,76,74,76,76,63,54),
(77,81,75,52,64,75,108,109,114,90,73,80,77,74,80,80,81,102,113,107,93,78,79,77,78,60,54,78,72,57,75,84,113,108,113,80,75,80,76,76,80,80,84,110,110,106,86,78,78,77,75,53,58,81,85,77,52,65,79,109,112,111,86,79,77,83,83,82,78,79,110,112,103,96,76,80,75,74,63,53),
(78,78,70,53,67,80,93,98,110,85,77,79,76,75,78,79,76,91,95,111,94,76,79,83,99,69,54,80,70,52,75,83,95,102,107,78,80,78,75,76,78,78,79,95,98,112,85,77,78,89,96,57,60,80,72,69,58,71,78,90,104,113,89,79,82,80,79,79,79,72,88,97,108,97,82,79,78,98,72,53),
(80,60,55,56,78,80,72,89,116,81,71,74,79,83,77,76,73,76,81,110,95,75,79,89,118,76,52,79,68,52,80,80,72,100,112,72,74,74,81,82,76,76,73,77,88,113,84,77,79,99,115,60,60,82,54,52,56,72,77,71,79,115,90,79,80,78,74,73,80,80,74,78,112,95,76,78,84,117,78,51),
(88,58,52,44,64,77,67,92,121,86,71,74,80,91,89,88,87,87,84,110,95,74,79,87,117,73,50,78,66,48,68,70,70,105,115,77,73,74,83,92,89,88,87,85,90,113,85,76,78,96,113,58,59,83,58,47,49,69,81,77,88,122,95,77,83,85,86,85,85,89,85,86,110,97,81,79,83,114,78,53),
(87,73,69,69,74,75,77,83,93,85,73,80,70,66,69,66,68,62,65,113,95,73,81,91,120,75,53,79,78,73,77,74,78,87,93,81,73,80,66,69,68,66,68,59,77,116,84,75,82,100,116,59,58,83,78,69,70,74,80,79,79,91,83,79,81,69,69,68,63,66,68,75,112,96,79,78,85,118,82,52),
(84,86,82,78,77,76,80,78,75,77,77,81,59,45,63,61,57,41,48,109,88,74,76,80,119,74,54,77,79,83,81,79,79,78,74,78,77,80,47,50,58,53,51,38,69,111,78,77,73,92,117,58,60,79,79,80,84,81,79,79,72,71,77,82,85,62,54,57,52,52,53,62,105,90,78,78,86,122,73,48),
(78,78,76,75,76,75,75,81,83,81,80,78,68,56,59,55,53,56,61,108,97,78,79,84,118,74,53,73,77,80,82,77,76,83,83,81,79,78,59,56,56,51,51,42,76,126,86,78,78,94,116,58,64,77,78,81,79,81,79,78,77,80,84,83,85,69,53,51,52,51,47,53,113,90,74,80,88,121,74,49),
(81,80,81,81,81,78,77,74,61,78,77,76,73,70,68,66,65,65,79,132,112,80,77,80,97,79,68,78,78,78,82,77,78,69,64,80,76,77,70,69,71,70,71,61,89,135,98,78,77,84,97,70,73,80,76,75,75,77,75,82,72,59,78,85,83,77,63,82,89,97,77,67,130,105,74,80,84,98,82,68),
(77,77,78,81,82,77,78,70,41,72,76,78,76,80,80,79,81,68,84,137,115,79,76,71,73,80,79,80,77,77,81,75,80,58,46,78,74,79,76,81,81,83,85,76,102,137,100,77,75,71,75,81,80,84,77,73,78,83,80,85,74,42,73,85,81,82,73,107,114,116,89,92,140,120,79,79,77,79,88,87),
(80,85,84,81,81,77,80,72,46,67,80,81,79,78,75,76,82,80,84,120,105,77,82,77,77,79,77,79,78,82,81,75,82,62,48,74,80,81,79,75,67,71,78,73,95,130,93,77,82,76,77,78,78,80,86,84,84,83,81,81,76,50,76,84,82,75,71,103,111,121,85,86,124,105,78,80,79,80,78,76),
(78,65,54,60,74,79,83,73,72,76,80,79,76,74,78,81,84,86,82,93,88,76,82,77,76,73,73,79,76,56,72,81,82,71,74,77,80,78,75,80,100,100,101,80,84,98,82,78,82,76,76,70,74,76,67,66,60,63,81,82,74,73,85,81,80,93,100,115,108,87,78,78,94,86,80,82,82,82,75,76));

CONSTANT SKY_R: my_background :=
((51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,51,50,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,48,51,56,48,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,50,50),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,50,51,45,42,54,54,50,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,53,51,51),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,52,50,67,74,53,53,50,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,51,51,52),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,47,55,44,176,244,101,41,55,50,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,47,38,48,46),
(51,51,51,51,51,51,51,51,51,51,51,51,53,49,50,70,39,80,246,255,210,42,45,57,51,50,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,43,78,162,81,61),
(51,51,51,51,51,51,51,51,51,51,51,51,52,45,169,230,67,168,232,175,239,201,73,30,51,52,50,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,53,42,163,255,178,174),
(51,51,51,51,51,51,51,51,51,51,51,52,45,63,238,255,208,241,200,205,197,255,193,125,63,49,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,48,194,255,247,248),
(51,51,51,51,51,51,51,51,51,51,51,52,48,72,240,251,248,244,247,233,159,189,252,255,151,42,54,50,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,52,54,35,194,255,249,252),
(51,51,51,51,51,51,51,51,51,51,49,53,40,94,249,253,250,251,251,241,249,245,249,255,219,60,48,56,55,53,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,50,47,49,43,126,240,255,251,248),
(51,51,51,51,51,51,51,51,51,51,54,46,93,234,251,254,247,249,249,253,254,255,250,250,226,45,49,38,50,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,50,52,59,44,90,249,254,252,254,254),
(51,51,51,51,51,51,51,51,51,51,58,42,176,255,250,251,255,255,253,252,254,251,253,255,227,145,218,129,42,51,49,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,50,55,49,48,29,121,255,248,255,248,233),
(51,51,51,51,51,51,51,51,51,48,44,35,195,255,248,255,215,200,254,254,254,255,231,197,241,248,255,242,71,35,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,44,84,116,165,255,248,255,214,169),
(51,51,51,51,51,51,51,52,45,64,176,196,237,251,251,235,189,194,161,188,246,254,217,189,216,255,247,255,170,91,49,52,50,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,53,43,78,232,255,254,254,253,247,206,253),
(51,51,51,51,51,51,51,53,44,165,255,253,242,248,255,234,234,246,199,231,247,252,249,254,180,238,253,253,255,234,73,48,53,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,54,38,144,255,249,201,197,250,245,246,255),
(51,51,51,51,51,51,51,51,49,217,255,230,166,188,221,251,252,247,250,252,255,253,255,235,170,194,255,252,241,255,125,42,55,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,55,34,169,255,222,192,195,154,239,255,253),
(51,51,51,51,51,51,52,49,60,227,255,198,234,186,191,253,252,249,250,248,251,251,252,248,251,241,250,253,249,255,172,38,54,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,51,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,53,41,187,255,233,243,227,217,253,246,255),
(51,51,51,51,51,51,52,46,73,245,255,252,253,239,255,255,255,255,255,255,255,255,255,255,255,255,255,255,252,255,174,41,53,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,55,52,51,54,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,45,199,255,252,254,254,255,255,254,255),
(51,51,51,51,51,51,52,46,73,199,201,201,200,204,204,206,206,209,209,209,209,210,211,211,211,212,214,214,212,223,127,47,55,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,51,57,43,38,49,48,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,46,79,92,90,91,93,92,93,93,94),
(51,51,51,51,51,51,51,51,48,49,44,41,42,44,45,43,43,45,46,45,45,47,47,48,49,48,48,48,47,51,50,44,50,51,51,51,51,51,51,51,51,51,51,51,51,51,53,51,51,45,151,166,50,53,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,50,54,49,43,41,41,43,43,43,43,42),
(51,51,51,51,51,51,51,51,51,49,52,54,53,52,56,55,55,53,52,52,52,51,51,51,52,52,51,51,51,51,47,53,49,51,51,51,51,51,51,51,51,51,51,51,51,50,44,55,43,77,247,255,123,26,57,53,50,51,51,51,51,51,51,51,51,51,51,51,51,51,48,51,52,54,55,56,56,55,55,53),
(51,51,51,51,51,51,51,51,51,51,50,50,50,50,50,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,38,102,215,72,158,226,202,239,120,32,44,49,53,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,53,44,182,255,211,232,208,197,220,240,146,87,49,57,50,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,50,54,35,181,255,253,247,252,208,169,228,255,209,59,53,52,50,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,53,51,54,47,73,218,254,243,245,253,246,248,247,244,250,74,27,53,55,46,49,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,54,52,57,209,255,249,252,253,249,252,253,248,251,246,97,97,62,49,57,48,50,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,49,48,29,81,255,249,252,242,239,255,254,253,252,240,246,206,255,184,39,49,58,49,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,53,48,61,107,144,253,247,250,190,183,208,215,255,243,171,208,255,248,247,101,41,50,53,51,51,51,51,51,51,50,51,53,51,51,50,51,51,51,51,51),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,54,45,166,255,251,250,255,238,226,234,175,223,253,248,254,197,233,255,251,255,159,38,53,51,51,51,53,49,51,54,54,46,53,49,55,51,51,51,51,51),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,62,231,255,209,184,218,247,252,249,250,255,255,250,250,192,189,249,254,255,235,67,48,52,51,51,50,54,50,48,49,58,48,59,50,51,51,51,51,51),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,53,44,77,249,240,208,208,175,245,248,249,249,251,251,251,246,241,228,244,253,249,254,100,41,53,51,51,52,51,51,26,129,254,73,40,53,50,51,51,51,51),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,53,40,89,255,253,253,249,249,255,255,255,255,255,255,255,255,255,255,255,255,254,255,98,41,53,51,51,51,52,171,120,185,221,208,74,43,53,50,51,51,51),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,53,44,78,174,173,175,177,173,175,176,175,175,176,178,176,175,175,176,176,177,180,176,68,48,52,47,51,43,71,247,244,236,203,211,234,136,44,55,50,48,49),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,53,48,33,37,37,37,38,38,38,38,38,39,40,40,40,40,40,40,40,39,36,51,52,50,53,58,40,104,249,252,253,245,226,255,232,46,44,53,49,51),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,52,51,51,51,51,51,51,51,51,51,51,51,51,52,51,51,51,51,51,51,54,57,52,52,52,52,52,52,52,52,52,52,52,52,52,52,52,52,53,54,48,50,51,51,43,54,225,254,255,255,254,254,255,233,128,98,46,53,53),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,53,48,49,51,52,50,51,51,51,51,51,51,51,52,55,45,53,51,51,50,52,48,45,52,54,53,52,52,52,52,52,52,52,52,52,52,52,52,52,52,51,50,57,52,51,51,56,118,254,249,220,213,231,254,220,221,255,236,73,39,52),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,46,50,58,56,45,50,50,53,51,51,51,50,47,52,44,41,89,45,53,50,52,50,53,54,52,52,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,52,49,56,205,246,246,245,227,204,202,251,242,203,237,251,225,83,44),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,31,185,187,41,53,54,48,51,51,51,52,55,42,82,113,216,122,40,63,49,51,51,50,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,53,41,93,254,211,187,221,255,249,248,249,249,209,221,244,255,162,39),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,51,50,183,159,209,230,156,50,45,54,50,52,51,52,57,40,148,255,224,242,142,29,58,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,54,38,112,255,245,245,250,255,255,255,255,255,255,255,252,255,176,34),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,48,58,232,255,237,198,242,213,52,46,54,49,50,53,36,56,225,245,241,255,221,113,44,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,46,78,142,138,140,142,140,142,144,145,145,145,150,143,147,101,45),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,53,57,40,138,251,252,254,252,255,247,93,54,55,48,52,46,70,192,246,225,220,238,216,247,121,40,50,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,47,39,39,39,38,38,38,38,38,37,38,38,38,40,46,51),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,44,59,223,255,232,234,249,246,224,235,190,44,55,55,37,124,255,228,255,255,255,242,255,205,46,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,54,54,54,54,54,54,54,54,54,54,54,54,53,52,51),
(51,51,51,51,51,51,51,51,51,51,51,51,51,53,42,108,224,240,248,218,203,231,249,208,239,255,170,50,51,49,68,120,117,115,122,117,121,120,103,50,50,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51),
(51,51,51,51,51,51,51,51,51,51,51,51,51,53,39,177,249,191,225,253,252,247,255,231,221,252,255,94,41,55,48,36,41,39,40,40,37,39,36,50,50,52,51,51,51,51,51,51,51,51,51,51,51,51,51,52,51,48,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51),
(51,51,51,51,51,51,51,51,51,51,51,51,51,52,44,193,253,237,242,255,252,254,255,255,255,253,255,111,39,53,52,55,54,54,53,53,54,54,53,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,50,53,59,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,50,79,92,93,91,91,87,89,89,90,91,96,91,59,49,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,53,51,47,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,42,41,44,41,43,43,44,44,42,38,40,46,48,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,50,51,47,49,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51),
(51,51,50,49,52,54,50,51,51,51,51,51,51,51,51,54,59,55,54,52,52,52,52,54,57,55,54,49,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,59,104,180,53,48,52,50,50,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51),
(51,51,52,50,50,54,52,51,51,51,51,51,51,51,51,51,50,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,56,34,146,238,220,186,54,49,53,49,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51),
(51,51,53,56,48,50,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,46,54,222,255,246,255,163,57,43,53,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51),
(51,52,49,56,57,48,56,50,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,51,51,51,51,51,51,51,52,48,62,179,246,224,234,227,239,184,54,50,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51),
(54,47,32,81,207,74,36,56,53,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,53,52,47,52,53,51,51,51,51,51,51,53,40,110,255,236,254,254,252,248,255,100,39,54,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51),
(38,111,144,154,242,199,65,42,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,49,58,53,49,50,51,51,51,51,51,51,52,48,69,103,105,110,108,110,110,109,69,48,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51),
(27,155,255,239,209,210,235,102,42,54,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,56,38,40,57,51,51,51,51,51,51,51,51,50,37,39,40,39,37,39,38,42,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51),
(65,206,255,248,247,239,255,168,30,52,53,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,50,53,44,112,102,40,54,51,50,51,51,51,51,51,50,54,54,55,54,52,53,56,56,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51),
(141,255,239,240,251,254,242,217,203,83,35,53,50,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,50,44,42,55,235,255,83,35,57,55,48,53,51,51,51,50,51,52,49,50,52,51,50,53,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51),
(215,255,228,200,221,254,219,216,255,200,78,49,54,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,50,53,191,119,124,229,216,216,84,34,49,56,52,51,51,51,51,51,51,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51),
(211,212,244,240,233,252,244,197,230,255,183,43,55,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,53,43,92,255,229,228,212,189,224,223,140,58,42,49,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,50,51,51,52,51,51,51,51,51),
(236,229,255,255,255,255,255,255,253,255,207,44,52,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,50,49,54,38,89,255,250,249,250,215,190,239,255,132,43,58,53,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,53,54,52,51,49,53,51,51,51,51),
(142,142,140,140,140,140,141,144,143,148,115,46,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,49,54,47,62,185,255,245,248,253,250,255,247,255,165,30,44,49,54,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,50,55,51,49,54,49,49,44,46,55,52,50),
(36,36,35,34,34,34,34,34,34,33,39,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,54,53,34,136,255,250,255,253,248,254,251,252,255,185,159,139,48,54,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,52,55,45,55,176,157,53,52,56,52),
(55,55,54,54,54,54,52,51,51,51,51,51,51,51,51,51,51,51,50,51,52,51,51,51,51,51,51,51,51,51,51,51,51,51,54,52,52,165,255,254,229,201,234,240,255,229,203,245,255,244,79,36,54,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,53,47,41,42,42,106,255,255,131,25,50,52),
(52,52,53,54,54,54,52,50,51,51,51,51,51,51,51,51,50,49,56,50,46,51,52,52,51,51,51,51,51,51,51,51,51,52,43,144,234,246,253,251,215,213,173,218,255,237,207,220,251,250,223,108,42,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,54,154,146,35,184,231,212,230,108,45,46),
(50,50,50,50,50,50,50,50,50,50,51,51,51,51,51,51,51,50,38,60,51,52,53,53,51,51,51,51,51,51,51,51,52,47,64,233,255,208,218,248,248,247,234,254,249,255,232,171,240,251,255,218,53,48,52,51,51,51,51,51,51,51,51,51,51,51,51,52,45,101,255,229,156,244,188,189,244,247,113,67),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,49,64,75,183,122,30,54,50,51,51,51,51,51,51,51,51,53,43,83,254,223,205,180,211,251,245,251,251,251,248,242,227,233,252,247,248,88,44,52,51,51,51,51,51,51,51,51,51,51,51,51,54,37,115,255,247,254,233,239,212,153,229,249,224),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,54,40,102,241,222,220,138,36,55,50,51,51,51,51,51,51,51,53,41,102,255,252,253,247,255,255,255,255,255,255,255,255,255,255,254,255,253,85,44,53,51,51,51,51,51,51,51,51,51,51,52,51,54,37,126,255,248,246,252,253,221,222,222,252,253),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,54,33,179,254,242,253,226,92,45,53,51,51,51,51,51,51,51,52,46,75,148,145,144,142,143,147,147,146,145,146,149,148,149,149,151,153,142,57,49,51,51,51,51,51,51,51,51,51,51,52,47,50,41,90,218,255,251,248,252,250,251,255,253,248,249),
(51,51,51,51,51,51,51,51,51,51,51,51,51,52,48,44,136,239,231,221,242,215,240,114,39,54,51,51,51,51,51,51,51,52,46,35,34,33,34,35,35,35,35,34,34,34,34,35,35,35,34,37,50,51,51,51,51,51,51,51,51,51,51,51,49,56,59,57,198,255,250,246,254,249,249,252,249,251,255,254),
(51,51,51,51,51,51,51,51,51,51,51,51,51,53,44,89,249,232,253,255,255,236,255,231,62,46,51,51,51,51,51,51,51,51,51,53,55,57,56,57,56,53,54,57,56,53,53,53,53,53,53,54,51,51,51,51,51,51,51,51,51,51,51,50,53,50,26,44,237,255,247,255,224,241,255,252,250,247,240,242),
(51,51,51,51,51,51,51,51,51,51,51,51,51,52,46,73,163,163,171,171,167,174,173,158,59,48,52,51,51,51,51,51,51,51,51,51,51,52,51,50,51,51,51,52,52,52,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,45,62,125,137,237,253,255,237,176,190,202,220,255,252,190,166),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,50,36,38,38,40,41,39,36,39,44,53,51,51,51,51,51,51,51,51,51,51,50,50,50,50,50,51,51,50,50,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,45,177,255,254,252,247,255,208,245,209,177,220,247,248,250,247),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,54,54,54,53,53,53,54,53,52,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,53,44,82,249,253,228,178,239,249,244,253,244,246,252,250,254,255,230),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,53,40,103,255,244,183,214,151,201,255,251,254,248,251,254,254,255,231),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,54,38,125,255,239,229,250,208,249,253,251,249,252,254,252,254,254,254),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,54,38,131,255,252,255,253,253,255,255,255,255,255,255,255,255,255,254),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,47,66,99,95,91,96,97,96,96,96,96,97,102,103,102,102,104),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,50,38,47,46,45,45,45,46,46,45,45,41,40,41,41,41),
(51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,52,50,50,49,50,51,51,50,51,51,51,52,52,52,52,53));

CONSTANT SKY_G: my_background :=
((190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,191,189,190,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,190,190),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,188,187,190,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,188,188,190),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,190,192,187,193,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,194,191,190),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,189,230,249,206,186,191,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,184,193,188),
(190,190,190,190,190,190,190,190,190,190,190,190,190,189,188,192,185,194,250,255,235,187,190,188,193,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,190,199,226,195,194),
(190,190,190,190,190,190,190,190,190,190,190,190,191,186,227,244,193,226,243,228,249,235,188,184,188,188,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,184,225,255,228,224),
(190,190,190,190,190,190,190,190,190,190,190,190,190,192,247,255,233,246,232,238,231,251,234,213,191,188,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,187,234,255,250,251),
(190,190,190,190,190,190,190,190,190,190,190,190,189,198,248,251,254,248,249,245,216,232,254,255,222,183,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,190,192,187,235,255,253,251),
(190,190,190,190,190,190,190,190,190,190,190,190,188,201,248,253,250,251,251,247,251,249,250,252,239,189,189,188,188,192,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,190,195,192,187,215,246,252,253,252),
(190,190,190,190,190,190,190,190,190,190,191,188,197,251,251,253,254,253,254,255,254,253,253,255,240,187,186,191,192,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,192,188,187,187,198,250,255,252,253,254),
(190,190,190,190,190,190,190,190,190,191,189,187,227,255,251,254,251,252,253,254,253,254,254,255,243,212,246,214,187,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,192,191,179,214,255,252,252,252,244),
(190,190,190,190,190,190,190,190,190,189,187,183,232,255,253,255,240,237,255,254,254,255,246,230,252,252,254,248,195,187,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,196,206,223,254,251,255,235,221),
(190,190,190,190,190,190,190,190,190,193,230,232,246,251,251,248,228,234,221,224,250,253,236,227,237,254,253,255,224,202,187,190,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,197,244,255,251,253,252,248,233,255),
(190,190,190,190,190,190,190,191,186,226,255,253,247,252,254,246,246,247,227,247,250,252,254,252,228,248,255,251,253,246,194,189,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,183,217,255,252,233,230,251,250,250,255),
(190,190,190,190,190,190,190,190,190,241,253,246,217,228,237,252,253,251,252,252,254,252,254,244,216,234,255,255,252,255,214,186,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,185,226,255,242,228,234,221,248,253,254),
(190,190,190,190,190,190,190,190,192,242,255,231,248,220,233,254,252,251,251,251,250,252,253,251,249,249,254,253,250,255,222,185,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,190,190,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,188,236,255,244,246,239,241,255,254,254),
(190,190,190,190,190,190,190,188,197,252,253,253,254,245,255,255,255,255,255,255,255,255,255,255,255,255,255,255,254,255,227,187,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,189,188,193,192,192,190,189,189,190,190,190,190,190,190,190,190,190,190,190,190,190,191,187,233,253,254,254,251,253,254,254,254),
(190,190,190,190,190,190,190,189,195,235,239,238,238,239,237,237,237,237,237,237,236,238,239,239,239,240,242,242,241,246,212,184,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,189,187,183,186,188,190,189,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,200,202,204,203,204,203,204,204,201),
(190,190,190,190,190,190,190,190,190,185,187,187,187,187,184,187,188,186,186,186,186,187,188,189,190,189,189,189,189,188,193,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,189,190,187,218,219,192,188,189,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,188,186,190,187,187,185,185,185,185,185),
(190,190,190,190,190,190,190,190,189,189,190,189,189,189,189,190,190,189,189,189,189,189,188,189,190,190,189,189,189,189,191,189,189,190,190,190,190,190,190,190,190,190,190,190,190,190,187,189,185,195,253,255,208,187,191,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,190,191,191,191,191,190,190,190),
(190,190,190,190,190,190,190,190,190,191,190,191,191,191,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,186,205,239,195,224,243,233,248,206,184,187,187,189,190,190,190,190,190,190,190,190,190,190,190,190,190,191,190,190,190,190,190,190,190,190),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,186,231,255,238,243,233,230,241,247,220,198,186,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,181,232,255,252,247,253,241,225,240,255,237,190,190,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,189,192,196,240,255,252,255,250,250,252,248,252,249,201,185,188,192,192,190,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,188,192,192,192,242,254,251,248,251,250,254,254,252,252,251,198,201,195,186,186,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,189,188,181,196,253,252,250,245,247,253,251,251,250,250,250,234,255,223,185,192,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,189,212,223,255,252,251,232,225,233,240,254,249,222,238,255,249,253,205,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,187,227,255,251,252,255,248,241,243,227,239,253,250,250,235,249,252,251,253,218,187,191,190,190,190,188,194,193,192,187,188,191,190,190,190,190,190,190,190),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,195,248,252,235,224,240,250,254,251,251,254,254,253,255,228,225,252,255,255,247,192,190,190,190,190,191,186,187,193,191,194,187,189,189,191,190,190,190,190),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,188,199,250,247,235,238,222,250,252,250,250,252,253,253,248,248,245,250,254,252,253,204,186,191,190,190,190,191,187,183,213,250,195,184,192,190,190,190,190,190),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,186,206,255,253,252,251,251,255,255,254,255,255,255,255,254,254,255,253,255,255,255,205,187,191,190,190,189,189,225,204,231,240,238,192,187,190,190,190,190,190),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,199,229,227,225,228,229,230,231,230,230,231,231,232,233,233,232,232,232,231,230,194,190,190,191,191,190,193,252,250,247,234,238,248,213,188,190,189,190,190),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,188,184,180,181,182,182,182,182,181,181,182,183,184,184,184,184,184,184,184,184,187,190,190,186,190,183,205,252,254,253,249,244,254,246,186,187,192,188,189),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,190,190,190,190,190,188,188,192,192,191,191,192,192,192,191,191,191,192,192,192,192,192,192,192,192,191,189,190,190,191,190,192,245,255,254,254,252,252,255,244,212,201,188,189,188),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,190,190,191,190,190,190,190,190,190,190,190,190,187,189,190,190,190,190,190,190,191,190,190,189,189,189,189,189,189,189,189,189,189,189,189,189,189,190,191,191,190,191,190,186,206,252,253,238,237,246,253,240,242,255,248,193,191,190),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,192,191,191,191,188,188,188,191,191,190,190,190,190,190,191,190,187,199,191,186,191,191,190,190,189,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,189,190,189,190,237,253,251,252,243,233,234,254,246,234,246,250,244,201,189),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,188,184,230,230,188,188,187,191,190,190,190,190,192,187,197,212,241,204,191,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,188,203,255,238,227,237,253,251,252,251,254,235,238,253,255,218,183),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,235,222,234,240,221,190,191,186,191,190,190,190,193,188,219,253,239,245,216,183,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,187,210,255,247,247,250,255,255,255,255,255,255,255,254,255,230,184),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,192,190,188,246,254,247,234,247,238,190,191,190,189,190,190,187,190,249,251,250,253,241,208,185,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,188,199,216,217,218,217,214,215,217,216,215,215,217,215,218,204,189),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,188,187,216,252,254,252,251,253,251,197,190,192,189,190,189,195,230,244,243,240,248,241,249,207,186,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,188,184,184,184,184,183,184,185,185,184,185,185,185,184,187,190),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,191,244,255,242,245,253,251,238,247,230,182,190,191,187,212,255,242,254,254,255,249,255,241,188,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,190),
(190,190,190,190,190,190,190,190,190,190,190,190,190,191,186,204,245,252,251,237,231,245,252,233,247,251,223,188,190,189,198,210,213,206,210,206,212,208,198,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,190),
(190,190,190,190,190,190,190,190,190,190,190,190,190,191,185,232,250,230,244,253,253,252,254,244,239,255,254,203,188,189,188,189,184,188,188,187,187,185,187,189,192,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,190,190,190,190,190,190,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,190),
(190,190,190,190,190,190,190,190,190,190,190,190,190,191,187,235,252,245,250,254,253,254,254,254,255,252,255,205,187,191,190,190,190,191,191,191,190,191,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,197,199,194,195,197,197,197,196,196,197,197,200,187,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,190,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,189,187,190,187,187,188,188,187,187,188,185,187,188,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,187,186,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190),
(190,190,189,191,189,189,189,190,190,190,190,190,190,190,190,188,190,191,188,190,192,191,191,191,191,191,190,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,190,193,204,227,184,190,191,191,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190),
(190,190,192,192,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,188,220,250,240,228,192,187,189,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190),
(190,190,194,191,185,190,186,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,189,242,252,250,252,221,189,191,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190),
(190,191,190,188,188,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,193,226,248,236,245,242,247,234,188,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190),
(190,190,186,201,241,194,188,190,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,190,191,188,190,190,190,190,190,190,190,191,186,207,254,247,255,254,252,250,255,201,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190),
(182,207,220,224,247,233,189,186,188,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,192,191,189,191,194,191,190,190,190,190,190,190,189,195,206,206,205,205,204,205,206,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190),
(185,219,255,246,239,235,244,207,191,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,192,193,187,186,189,190,190,190,190,190,190,191,186,187,186,187,186,184,183,186,190,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190),
(189,236,252,252,250,247,255,225,182,191,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,192,189,186,202,203,190,191,190,190,190,190,190,190,190,192,190,192,189,191,194,195,189,189,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190),
(214,255,247,245,253,253,248,237,239,196,186,189,188,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,189,188,187,185,192,242,254,195,189,194,190,191,190,190,190,190,190,188,191,189,189,190,190,189,188,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190),
(243,252,242,230,238,254,235,238,251,238,195,187,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,189,187,230,210,211,243,240,241,194,182,189,187,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190),
(232,234,248,251,247,253,250,232,245,255,230,186,192,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,186,200,255,245,244,236,232,244,240,212,192,190,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190),
(248,247,254,253,255,255,254,251,252,255,241,186,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,190,189,186,200,251,251,249,255,238,228,250,255,215,185,193,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,188,190,190,191,192,190,191,191,190),
(217,217,218,218,217,218,217,217,217,219,209,188,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,192,186,191,230,253,252,252,250,251,254,251,255,221,180,189,191,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,188,190,192,188,192,185,184,191,188,190,188),
(187,187,185,185,185,185,185,185,185,184,186,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,192,192,186,217,255,254,252,253,252,254,252,249,255,226,221,211,184,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,187,193,189,189,190,190,226,220,187,189,187,188),
(192,192,190,190,190,190,190,191,191,191,190,190,190,190,190,190,190,190,190,190,190,191,190,190,190,190,190,190,190,190,190,190,190,190,188,187,186,222,253,254,245,230,246,249,254,244,233,249,254,254,197,185,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,188,181,186,186,206,254,255,208,181,192,191),
(188,188,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,189,191,188,191,190,190,190,190,190,190,190,190,190,190,191,186,216,246,251,253,252,237,238,222,235,254,243,238,242,252,248,243,206,187,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,191,222,217,185,233,242,241,246,204,186,189),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,190,186,191,191,191,190,190,190,190,190,190,190,190,190,189,193,247,253,233,240,251,249,251,247,255,254,255,246,222,248,255,255,242,188,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,187,203,255,245,220,252,226,227,245,250,203,193),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,193,191,230,207,186,191,188,190,190,190,190,190,190,190,190,190,188,199,249,243,234,223,236,253,251,253,251,251,252,249,245,244,252,252,251,199,187,191,190,190,190,190,190,190,190,190,190,190,190,190,191,187,212,253,251,251,246,248,238,218,244,251,244),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,186,205,248,239,244,212,185,190,190,190,190,190,190,190,190,190,191,187,206,255,254,253,248,255,255,255,254,255,255,255,255,254,255,255,255,255,200,187,191,190,190,190,190,190,190,190,190,190,190,190,190,192,180,210,255,251,253,250,255,240,238,245,254,253),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,184,225,255,250,251,240,201,186,189,191,190,190,190,190,190,190,190,188,195,220,217,215,220,217,218,221,222,221,220,221,219,221,219,224,224,220,191,190,190,190,190,190,190,190,190,190,190,190,189,189,187,189,202,242,253,251,250,252,249,250,251,251,252,251),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,190,209,250,242,237,250,240,251,203,184,190,190,190,190,190,190,190,190,190,187,182,182,181,181,182,182,182,182,182,182,182,182,183,183,183,183,185,190,190,190,190,190,190,190,190,190,190,190,190,188,190,190,192,239,255,252,253,250,252,248,252,253,249,251,253),
(190,190,190,190,190,190,190,190,190,190,190,190,190,191,186,198,255,247,254,251,255,244,255,244,189,190,190,190,190,190,190,190,190,190,189,189,191,192,192,193,191,189,190,193,193,190,190,190,190,190,190,191,190,190,190,190,190,190,190,190,190,190,190,190,191,192,187,192,247,254,253,250,245,247,254,252,252,253,249,246),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,199,221,220,220,223,225,227,227,220,191,189,190,190,190,190,190,190,190,190,189,189,189,190,189,188,189,189,189,191,191,191,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,188,190,206,215,248,253,253,242,222,228,232,240,252,249,229,225),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,187,184,187,185,185,184,186,184,184,189,189,190,190,190,190,190,190,190,190,190,190,189,189,189,188,189,190,190,189,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,230,255,252,253,252,253,237,248,239,224,236,253,253,251,249),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,191,191,191,191,191,191,191,191,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,188,198,252,251,239,221,241,252,252,253,250,250,253,254,255,255,246),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,187,208,253,249,226,241,218,235,255,253,251,251,254,255,255,255,244),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,185,212,255,246,244,250,237,247,253,252,251,252,255,252,255,255,253),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,185,215,255,253,254,253,253,255,255,255,254,254,255,254,255,255,255),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,192,196,198,199,201,204,203,203,203,203,203,202,202,201,201,202),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,185,187,188,187,186,186,186,187,186,186,186,187,187,187,187,188),
(190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,192,191,188,188,189,190,190,189,190,190,190,189,189,189,189,190));

CONSTANT SKY_B: my_background :=
((247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,246,245,245,248,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,249,248),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,245,250,250,247,249,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,246,247),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,246,245,245,240,249,246,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,251,245,245),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,248,247,244,249,240,249,247,247,247,246,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,243,252,247),
(247,247,247,247,247,247,247,247,247,247,247,247,247,248,246,242,250,241,248,253,244,235,250,249,246,250,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,246,245,246,238,243),
(247,247,247,247,247,247,247,247,247,247,247,246,249,242,243,244,240,245,247,233,245,246,240,248,248,245,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,245,250,254,245,242),
(247,247,247,247,247,247,247,247,247,247,247,247,249,240,243,244,242,245,243,244,240,251,244,235,243,249,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,248,247,251,250,251),
(247,247,247,247,247,247,247,247,247,247,247,247,248,247,251,252,251,248,250,243,227,240,250,250,242,246,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,244,243,252,250,253),
(247,247,247,247,247,247,247,247,247,247,246,247,248,238,244,247,253,251,251,248,253,247,246,247,243,242,252,246,248,249,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,247,247,247,244,241,248,249,254,251),
(247,247,247,247,247,247,247,247,247,247,249,251,238,246,252,254,249,248,252,253,254,254,255,250,250,244,242,249,252,246,248,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,250,250,250,245,252,252,249,249,253),
(247,247,247,247,247,247,247,247,247,247,250,249,247,253,252,251,251,252,253,254,254,250,250,253,242,240,247,238,243,247,248,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,251,247,249,242,249,252,252,248,245),
(247,247,247,247,247,247,247,247,247,247,246,244,243,252,253,250,247,245,254,254,255,251,246,243,248,248,248,245,242,249,246,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,244,246,237,245,246,252,251,254,242,239),
(247,247,247,247,247,247,247,247,249,245,244,249,246,248,254,249,233,239,233,239,250,251,240,234,242,251,254,255,239,235,245,248,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,245,241,251,247,249,250,249,250,235,255),
(247,247,247,247,247,247,247,248,242,241,247,240,251,252,249,248,247,250,236,251,249,250,255,250,235,250,254,251,250,248,241,251,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,245,247,253,253,238,240,251,251,252,255),
(247,247,247,247,247,247,247,248,245,243,253,247,227,238,243,249,251,251,248,245,254,252,252,245,235,238,255,254,251,252,242,251,248,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,241,252,245,231,240,233,249,254,254),
(247,247,247,247,247,247,247,247,245,244,252,238,249,234,241,252,250,253,249,247,252,249,246,251,247,246,253,252,252,252,243,251,248,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,246,246,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,249,246,248,244,246,254,250,255),
(247,247,247,247,247,247,247,247,242,249,248,250,249,242,255,253,253,253,253,254,253,252,251,252,249,250,252,251,250,251,242,248,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,250,251,250,249,250,248,251,251,249,247,247,247,247,247,247,247,247,247,247,247,247,247,247,246,247,248,248,246,242,245,244,244,248),
(247,247,247,247,247,247,247,247,242,246,247,250,250,250,248,245,246,246,246,246,246,248,249,248,248,249,251,250,250,252,246,248,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,250,251,245,244,245,253,250,251,250,247,247,247,247,247,247,247,247,247,247,247,247,247,248,244,240,239,247,246,243,243,243,243,248),
(247,247,247,247,247,247,247,247,248,244,243,245,245,242,241,243,244,244,244,244,244,245,245,245,245,245,244,244,244,243,247,250,246,247,247,247,247,247,247,247,247,247,247,247,247,247,247,252,252,248,241,242,241,249,251,250,247,247,247,247,247,247,247,247,247,247,247,247,247,247,245,250,251,242,243,250,250,250,250,247),
(247,247,247,247,247,247,247,247,244,250,251,250,250,248,251,250,250,249,249,249,249,249,249,248,248,248,247,248,247,248,250,251,247,247,247,247,247,247,247,247,247,247,247,247,247,245,246,244,252,247,246,253,239,247,254,248,245,248,247,247,247,247,247,247,247,247,247,247,247,247,248,247,248,252,251,249,249,248,248,250),
(247,247,247,247,247,247,247,247,246,246,246,246,246,246,246,247,248,248,248,248,248,247,247,247,247,248,248,248,248,248,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,243,245,242,239,244,246,242,244,238,241,248,245,252,247,247,247,247,247,247,247,247,247,247,247,247,247,247,246,247,247,247,247,246,246,247),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,247,242,248,243,247,240,240,245,239,240,240,250,251,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,246,247,250,252,253,250,251,240,237,243,252,240,248,246,248,246,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,247,246,246,249,243,246,251,246,250,248,251,242,244,253,250,248,248,247,250,247,246,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,249,249,250,244,242,247,252,253,250,254,252,251,253,247,249,247,238,237,250,245,248,248,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,245,251,249,251,242,253,253,252,250,247,253,249,252,253,249,250,244,254,243,239,253,251,246,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,246,251,241,244,242,253,253,253,229,226,241,245,252,249,226,239,250,252,243,230,237,251,247,247,247,247,247,247,247,247,246,246,247,247,247,247,247,247,247,247),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,245,246,250,250,250,249,249,241,247,228,244,251,248,251,243,247,250,255,251,240,244,247,247,247,247,247,248,245,248,252,251,248,249,249,247,247,247,247,247),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,245,249,249,238,237,244,250,254,250,251,253,255,253,248,239,236,251,255,254,249,244,248,247,247,247,249,246,248,251,241,232,246,243,249,248,247,247,247,247),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,248,251,247,236,243,237,249,252,251,251,254,254,254,250,246,247,250,254,254,251,246,248,247,247,247,250,248,247,248,245,250,236,249,246,246,247,247,247,247),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,249,245,245,250,250,247,244,250,250,249,246,254,254,254,253,245,246,247,254,253,252,246,247,247,247,246,250,243,240,237,241,235,246,237,247,247,247,247,247,247),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,249,245,242,251,249,246,249,249,248,249,248,250,251,249,248,249,248,248,249,246,240,246,248,247,247,244,243,251,246,250,248,240,241,249,243,246,251,249,245,246),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,250,247,245,246,247,246,246,246,249,250,250,251,249,247,247,247,247,248,247,242,243,246,247,245,252,243,238,250,251,251,252,248,249,247,240,251,250,250,247),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,250,252,246,246,246,249,249,249,249,248,247,247,247,247,247,247,247,247,247,246,247,247,247,247,247,249,243,249,253,255,254,254,251,253,248,243,245,247,253,249),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,246,246,248,249,246,248,248,247,247,247,247,247,247,247,247,248,247,247,247,247,247,247,246,244,246,249,249,247,247,247,247,248,248,248,248,249,249,249,249,249,249,248,245,252,248,247,250,240,240,246,248,244,244,246,251,245,247,252,249,240,248,249),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,249,248,247,247,242,246,246,247,249,247,247,247,248,249,248,252,246,245,242,251,250,247,247,246,248,249,248,248,248,248,248,248,247,247,247,247,247,247,247,247,247,247,247,249,247,247,249,239,247,249,246,248,242,237,236,248,244,239,250,250,244,242,244),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,243,242,244,241,247,247,241,247,247,247,247,248,246,250,247,239,242,240,244,250,242,248,247,247,246,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,240,236,245,255,253,250,249,252,238,243,252,248,248,247),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,250,244,241,242,240,242,245,252,252,247,247,247,246,247,251,244,249,245,249,241,244,253,246,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,243,249,245,241,245,250,249,252,252,250,252,249,249,252,241,245),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,244,238,246,253,247,238,247,241,248,244,246,248,247,247,250,239,247,242,249,250,239,237,243,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,245,240,241,246,244,241,242,242,239,244,245,241,243,238,240,247),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,247,247,242,252,253,250,251,254,247,235,241,252,246,247,246,238,243,246,245,245,251,245,251,238,242,246,248,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,251,249,249,250,249,249,249,249,249,250,251,250,250,248,252,249),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,246,246,248,249,251,243,245,251,252,245,243,245,242,247,246,246,244,249,239,252,249,245,244,243,241,247,249,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,250,252,251,251,251,251,251,251,251,251,251,251,251,252,251,248),
(247,247,247,247,247,247,247,247,247,247,247,247,247,248,245,244,249,251,249,239,238,246,251,243,247,247,241,246,247,248,241,236,243,239,246,245,241,246,240,246,248,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,250,251,251,251,251,251,251,251,251,251,251,251,251,251,251,248),
(247,247,247,247,247,247,247,247,247,247,247,247,247,248,245,247,243,239,248,252,253,252,254,246,246,254,248,243,248,245,246,250,245,251,250,250,250,250,246,248,246,248,247,247,247,247,247,247,247,247,247,247,247,247,247,246,249,249,247,247,247,247,247,247,249,250,250,250,250,250,250,250,250,250,250,250,250,250,250,248),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,245,243,245,242,249,250,249,250,249,249,249,247,246,242,246,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,249,249,245,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,239,241,244,243,241,240,240,240,241,242,244,240,246,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,249,245,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,245,244,250,247,250,249,249,249,248,247,247,245,245,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,250,250,245,248,248,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247),
(247,247,246,247,246,248,247,247,247,247,247,247,247,247,247,248,247,248,247,250,250,250,250,250,250,250,249,246,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,246,241,240,240,241,244,243,248,246,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247),
(247,247,248,248,249,253,249,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,246,247,238,249,241,242,247,248,249,248,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247),
(247,247,250,248,247,252,245,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,239,246,251,251,249,241,242,248,244,248,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247),
(247,248,246,249,244,248,251,246,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,246,239,249,244,243,248,241,244,239,246,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247),
(249,249,246,244,249,243,250,249,249,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,249,250,250,250,248,247,247,247,247,247,247,247,247,240,250,247,249,251,249,246,252,237,248,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247),
(241,247,245,241,241,243,240,253,242,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,246,246,245,246,252,248,247,247,247,247,247,247,247,247,240,245,251,249,249,248,236,245,249,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247),
(250,247,243,247,238,241,246,245,245,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,246,248,255,248,251,245,246,247,247,247,247,247,247,247,250,248,249,249,249,246,247,248,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247),
(242,246,250,251,249,249,249,243,244,248,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,248,247,238,236,246,248,246,246,247,247,247,247,247,246,247,246,244,244,245,246,250,251,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247),
(243,251,247,247,252,249,247,242,248,241,247,249,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,249,251,249,240,238,243,249,245,241,248,246,246,251,249,247,247,247,247,247,249,249,249,249,248,247,248,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247),
(246,248,242,237,242,255,238,243,249,245,242,250,251,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,249,253,245,246,240,243,241,247,247,236,249,251,244,249,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247),
(233,243,246,250,247,254,253,233,247,250,240,248,252,246,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,249,251,250,245,245,248,238,234,244,246,239,243,245,247,248,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247),
(244,244,252,252,250,247,248,251,250,252,249,246,249,246,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,245,247,251,254,239,245,253,252,248,236,237,247,252,243,252,246,245,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,247,247,248,246,247,249,247,246,247,248,247),
(243,243,244,243,247,249,245,243,243,243,245,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,246,245,242,243,254,252,249,252,254,254,254,249,242,242,248,249,249,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,249,246,247,249,250,245,244,247,247,250,250),
(248,248,246,246,245,245,246,246,246,246,246,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,253,250,246,242,250,252,251,251,251,250,253,253,255,241,241,243,245,246,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,246,255,250,245,251,247,240,246,248,254,251,250),
(252,252,251,250,251,251,250,250,250,250,249,247,247,247,247,247,247,247,247,248,246,247,247,247,247,247,247,247,247,247,247,247,247,247,245,250,241,242,254,252,249,238,244,249,254,244,235,249,249,247,237,246,248,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,249,247,241,245,245,241,251,240,241,242,248,251),
(248,248,249,249,249,249,249,249,249,249,248,247,247,247,247,247,247,246,245,244,250,246,248,247,247,247,247,247,247,247,247,247,247,248,244,244,247,249,250,251,240,243,233,242,253,240,239,244,251,247,246,243,246,248,247,247,247,247,247,247,247,247,247,247,247,247,247,246,250,246,245,239,245,246,245,243,247,238,247,253),
(246,246,246,246,247,248,247,246,246,246,247,247,247,247,247,247,248,244,249,248,240,250,252,247,247,247,247,247,247,247,247,247,247,247,246,248,252,237,242,252,252,249,245,255,253,250,247,232,248,250,254,247,243,249,247,247,247,247,247,247,247,247,247,247,247,247,247,247,246,249,249,248,241,250,232,239,248,250,237,239),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,244,238,244,247,248,245,248,247,247,247,247,247,247,247,247,247,247,242,252,244,236,231,240,250,249,252,251,251,252,251,247,247,255,253,250,243,246,247,247,247,247,247,247,247,247,247,247,247,247,247,247,246,243,246,248,248,246,246,244,233,245,246,252),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,244,245,239,247,239,247,247,248,247,247,247,247,247,247,247,247,248,245,251,251,251,248,252,250,254,253,254,255,251,248,251,253,254,254,251,242,246,247,247,247,247,247,247,247,247,247,247,247,247,246,248,243,238,255,253,249,253,251,240,246,247,250,252),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,245,247,241,241,249,251,245,248,245,247,245,244,248,247,247,247,247,247,247,248,244,245,248,246,247,246,249,247,248,244,246,248,245,250,248,247,246,245,244,249,247,247,247,247,247,247,247,247,247,247,246,248,249,248,239,248,249,249,250,254,251,253,250,250,251,251),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,239,251,246,241,253,238,244,240,247,250,247,247,247,247,247,247,247,247,249,250,248,247,248,249,248,249,248,243,243,243,244,244,245,245,245,246,247,247,247,247,247,247,247,247,247,247,247,247,249,245,246,244,244,253,249,252,251,246,253,251,250,249,253,254),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,242,247,235,249,248,250,244,247,249,245,250,246,247,247,247,247,247,247,247,249,250,252,253,253,253,252,250,250,249,249,246,246,246,246,246,246,247,247,247,247,247,247,247,247,247,247,247,247,247,248,251,248,242,249,255,251,254,245,250,252,246,250,253,251,249),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,246,243,246,246,246,244,250,250,245,248,245,247,247,247,247,247,247,247,247,250,251,252,252,251,251,251,252,251,247,248,248,248,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,243,243,245,245,252,255,245,227,239,242,245,252,254,230,230),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,249,243,246,245,244,241,245,248,246,249,249,247,247,247,247,247,247,247,247,248,249,248,248,247,247,248,249,248,246,246,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,247,240,253,252,245,251,252,239,251,242,235,239,252,253,253,251),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,247,247,248,248,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,244,250,242,242,240,246,249,253,250,251,248,250,253,255,255,248),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,243,247,250,231,243,231,236,251,248,251,248,254,255,255,255,246),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,248,248,245,248,244,247,252,252,252,252,255,252,255,255,248),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,245,248,252,251,249,251,250,251,250,250,251,250,252,252,249),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,246,237,238,241,242,244,243,243,244,245,245,246,246,246,246,247),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,252,250,251,250,249,250,251,251,252,251,249,249,249,249,249),
(247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,247,248,245,247,244,245,246,246,247,247,248,247,246,246,246,246,247));

END background;